magic
tech sky130A
magscale 1 2
timestamp 1755619384
<< viali >>
rect 18245 10013 18279 10047
rect 18429 9877 18463 9911
rect 10701 3621 10735 3655
rect 10241 3553 10275 3587
rect 10333 3485 10367 3519
rect 10241 3145 10275 3179
rect 9873 3009 9907 3043
rect 10333 3009 10367 3043
rect 10425 3009 10459 3043
rect 10701 3009 10735 3043
rect 10885 3009 10919 3043
rect 9965 2941 9999 2975
rect 10609 2941 10643 2975
rect 10793 2941 10827 2975
rect 10517 2805 10551 2839
rect 9321 2601 9355 2635
rect 10149 2601 10183 2635
rect 11069 2601 11103 2635
rect 9965 2533 9999 2567
rect 9137 2397 9171 2431
rect 9781 2397 9815 2431
rect 10057 2397 10091 2431
rect 10701 2397 10735 2431
rect 11253 2397 11287 2431
rect 10517 2261 10551 2295
<< metal1 >>
rect 1104 17434 18860 17456
rect 1104 17382 3610 17434
rect 3662 17382 3674 17434
rect 3726 17382 3738 17434
rect 3790 17382 3802 17434
rect 3854 17382 3866 17434
rect 3918 17382 13610 17434
rect 13662 17382 13674 17434
rect 13726 17382 13738 17434
rect 13790 17382 13802 17434
rect 13854 17382 13866 17434
rect 13918 17382 18860 17434
rect 1104 17360 18860 17382
rect 1104 16890 18860 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 18860 16890
rect 1104 16816 18860 16838
rect 1104 16346 18860 16368
rect 1104 16294 3610 16346
rect 3662 16294 3674 16346
rect 3726 16294 3738 16346
rect 3790 16294 3802 16346
rect 3854 16294 3866 16346
rect 3918 16294 13610 16346
rect 13662 16294 13674 16346
rect 13726 16294 13738 16346
rect 13790 16294 13802 16346
rect 13854 16294 13866 16346
rect 13918 16294 18860 16346
rect 1104 16272 18860 16294
rect 1104 15802 18860 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 18860 15802
rect 1104 15728 18860 15750
rect 1104 15258 18860 15280
rect 1104 15206 3610 15258
rect 3662 15206 3674 15258
rect 3726 15206 3738 15258
rect 3790 15206 3802 15258
rect 3854 15206 3866 15258
rect 3918 15206 13610 15258
rect 13662 15206 13674 15258
rect 13726 15206 13738 15258
rect 13790 15206 13802 15258
rect 13854 15206 13866 15258
rect 13918 15206 18860 15258
rect 1104 15184 18860 15206
rect 1104 14714 18860 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 18860 14714
rect 1104 14640 18860 14662
rect 1104 14170 18860 14192
rect 1104 14118 3610 14170
rect 3662 14118 3674 14170
rect 3726 14118 3738 14170
rect 3790 14118 3802 14170
rect 3854 14118 3866 14170
rect 3918 14118 13610 14170
rect 13662 14118 13674 14170
rect 13726 14118 13738 14170
rect 13790 14118 13802 14170
rect 13854 14118 13866 14170
rect 13918 14118 18860 14170
rect 1104 14096 18860 14118
rect 1104 13626 18860 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 18860 13626
rect 1104 13552 18860 13574
rect 1104 13082 18860 13104
rect 1104 13030 3610 13082
rect 3662 13030 3674 13082
rect 3726 13030 3738 13082
rect 3790 13030 3802 13082
rect 3854 13030 3866 13082
rect 3918 13030 13610 13082
rect 13662 13030 13674 13082
rect 13726 13030 13738 13082
rect 13790 13030 13802 13082
rect 13854 13030 13866 13082
rect 13918 13030 18860 13082
rect 1104 13008 18860 13030
rect 1104 12538 18860 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 18860 12538
rect 1104 12464 18860 12486
rect 1104 11994 18860 12016
rect 1104 11942 3610 11994
rect 3662 11942 3674 11994
rect 3726 11942 3738 11994
rect 3790 11942 3802 11994
rect 3854 11942 3866 11994
rect 3918 11942 13610 11994
rect 13662 11942 13674 11994
rect 13726 11942 13738 11994
rect 13790 11942 13802 11994
rect 13854 11942 13866 11994
rect 13918 11942 18860 11994
rect 1104 11920 18860 11942
rect 1104 11450 18860 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 18860 11450
rect 1104 11376 18860 11398
rect 1104 10906 18860 10928
rect 1104 10854 3610 10906
rect 3662 10854 3674 10906
rect 3726 10854 3738 10906
rect 3790 10854 3802 10906
rect 3854 10854 3866 10906
rect 3918 10854 13610 10906
rect 13662 10854 13674 10906
rect 13726 10854 13738 10906
rect 13790 10854 13802 10906
rect 13854 10854 13866 10906
rect 13918 10854 18860 10906
rect 1104 10832 18860 10854
rect 1104 10362 18860 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 18860 10362
rect 1104 10288 18860 10310
rect 10686 10004 10692 10056
rect 10744 10044 10750 10056
rect 18233 10047 18291 10053
rect 18233 10044 18245 10047
rect 10744 10016 18245 10044
rect 10744 10004 10750 10016
rect 18233 10013 18245 10016
rect 18279 10013 18291 10047
rect 18233 10007 18291 10013
rect 18414 9868 18420 9920
rect 18472 9868 18478 9920
rect 1104 9818 18860 9840
rect 1104 9766 3610 9818
rect 3662 9766 3674 9818
rect 3726 9766 3738 9818
rect 3790 9766 3802 9818
rect 3854 9766 3866 9818
rect 3918 9766 13610 9818
rect 13662 9766 13674 9818
rect 13726 9766 13738 9818
rect 13790 9766 13802 9818
rect 13854 9766 13866 9818
rect 13918 9766 18860 9818
rect 1104 9744 18860 9766
rect 1104 9274 18860 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 18860 9274
rect 1104 9200 18860 9222
rect 1104 8730 18860 8752
rect 1104 8678 3610 8730
rect 3662 8678 3674 8730
rect 3726 8678 3738 8730
rect 3790 8678 3802 8730
rect 3854 8678 3866 8730
rect 3918 8678 13610 8730
rect 13662 8678 13674 8730
rect 13726 8678 13738 8730
rect 13790 8678 13802 8730
rect 13854 8678 13866 8730
rect 13918 8678 18860 8730
rect 1104 8656 18860 8678
rect 1104 8186 18860 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 18860 8186
rect 1104 8112 18860 8134
rect 1104 7642 18860 7664
rect 1104 7590 3610 7642
rect 3662 7590 3674 7642
rect 3726 7590 3738 7642
rect 3790 7590 3802 7642
rect 3854 7590 3866 7642
rect 3918 7590 13610 7642
rect 13662 7590 13674 7642
rect 13726 7590 13738 7642
rect 13790 7590 13802 7642
rect 13854 7590 13866 7642
rect 13918 7590 18860 7642
rect 1104 7568 18860 7590
rect 1104 7098 18860 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 18860 7098
rect 1104 7024 18860 7046
rect 1104 6554 18860 6576
rect 1104 6502 3610 6554
rect 3662 6502 3674 6554
rect 3726 6502 3738 6554
rect 3790 6502 3802 6554
rect 3854 6502 3866 6554
rect 3918 6502 13610 6554
rect 13662 6502 13674 6554
rect 13726 6502 13738 6554
rect 13790 6502 13802 6554
rect 13854 6502 13866 6554
rect 13918 6502 18860 6554
rect 1104 6480 18860 6502
rect 1104 6010 18860 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 18860 6010
rect 1104 5936 18860 5958
rect 1104 5466 18860 5488
rect 1104 5414 3610 5466
rect 3662 5414 3674 5466
rect 3726 5414 3738 5466
rect 3790 5414 3802 5466
rect 3854 5414 3866 5466
rect 3918 5414 13610 5466
rect 13662 5414 13674 5466
rect 13726 5414 13738 5466
rect 13790 5414 13802 5466
rect 13854 5414 13866 5466
rect 13918 5414 18860 5466
rect 1104 5392 18860 5414
rect 1104 4922 18860 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 18860 4922
rect 1104 4848 18860 4870
rect 1104 4378 18860 4400
rect 1104 4326 3610 4378
rect 3662 4326 3674 4378
rect 3726 4326 3738 4378
rect 3790 4326 3802 4378
rect 3854 4326 3866 4378
rect 3918 4326 13610 4378
rect 13662 4326 13674 4378
rect 13726 4326 13738 4378
rect 13790 4326 13802 4378
rect 13854 4326 13866 4378
rect 13918 4326 18860 4378
rect 1104 4304 18860 4326
rect 1104 3834 18860 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 18860 3834
rect 1104 3760 18860 3782
rect 10686 3612 10692 3664
rect 10744 3612 10750 3664
rect 10226 3544 10232 3596
rect 10284 3544 10290 3596
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 10321 3519 10379 3525
rect 10321 3516 10333 3519
rect 10100 3488 10333 3516
rect 10100 3476 10106 3488
rect 10321 3485 10333 3488
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 1104 3290 18860 3312
rect 1104 3238 3610 3290
rect 3662 3238 3674 3290
rect 3726 3238 3738 3290
rect 3790 3238 3802 3290
rect 3854 3238 3866 3290
rect 3918 3238 13610 3290
rect 13662 3238 13674 3290
rect 13726 3238 13738 3290
rect 13790 3238 13802 3290
rect 13854 3238 13866 3290
rect 13918 3238 18860 3290
rect 1104 3216 18860 3238
rect 10226 3136 10232 3188
rect 10284 3176 10290 3188
rect 10284 3148 10456 3176
rect 10284 3136 10290 3148
rect 9861 3043 9919 3049
rect 9861 3009 9873 3043
rect 9907 3009 9919 3043
rect 9861 3003 9919 3009
rect 9876 2904 9904 3003
rect 10318 3000 10324 3052
rect 10376 3000 10382 3052
rect 10428 3049 10456 3148
rect 10413 3043 10471 3049
rect 10413 3009 10425 3043
rect 10459 3009 10471 3043
rect 10689 3043 10747 3049
rect 10689 3040 10701 3043
rect 10413 3003 10471 3009
rect 10520 3012 10701 3040
rect 9950 2932 9956 2984
rect 10008 2972 10014 2984
rect 10520 2972 10548 3012
rect 10689 3009 10701 3012
rect 10735 3009 10747 3043
rect 10689 3003 10747 3009
rect 10873 3043 10931 3049
rect 10873 3009 10885 3043
rect 10919 3009 10931 3043
rect 10873 3003 10931 3009
rect 10008 2944 10548 2972
rect 10597 2975 10655 2981
rect 10008 2932 10014 2944
rect 10597 2941 10609 2975
rect 10643 2972 10655 2975
rect 10781 2975 10839 2981
rect 10781 2972 10793 2975
rect 10643 2944 10793 2972
rect 10643 2941 10655 2944
rect 10597 2935 10655 2941
rect 10781 2941 10793 2944
rect 10827 2941 10839 2975
rect 10781 2935 10839 2941
rect 10888 2904 10916 3003
rect 11054 2904 11060 2916
rect 9876 2876 11060 2904
rect 11054 2864 11060 2876
rect 11112 2864 11118 2916
rect 10505 2839 10563 2845
rect 10505 2805 10517 2839
rect 10551 2836 10563 2839
rect 10686 2836 10692 2848
rect 10551 2808 10692 2836
rect 10551 2805 10563 2808
rect 10505 2799 10563 2805
rect 10686 2796 10692 2808
rect 10744 2796 10750 2848
rect 1104 2746 18860 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 18860 2746
rect 1104 2672 18860 2694
rect 9309 2635 9367 2641
rect 9309 2601 9321 2635
rect 9355 2632 9367 2635
rect 10042 2632 10048 2644
rect 9355 2604 10048 2632
rect 9355 2601 9367 2604
rect 9309 2595 9367 2601
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 10137 2635 10195 2641
rect 10137 2601 10149 2635
rect 10183 2632 10195 2635
rect 10318 2632 10324 2644
rect 10183 2604 10324 2632
rect 10183 2601 10195 2604
rect 10137 2595 10195 2601
rect 10318 2592 10324 2604
rect 10376 2592 10382 2644
rect 11054 2592 11060 2644
rect 11112 2592 11118 2644
rect 9950 2524 9956 2576
rect 10008 2524 10014 2576
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 9088 2400 9137 2428
rect 9088 2388 9094 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9732 2400 9781 2428
rect 9732 2388 9738 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 10042 2388 10048 2440
rect 10100 2388 10106 2440
rect 10686 2388 10692 2440
rect 10744 2388 10750 2440
rect 10962 2388 10968 2440
rect 11020 2428 11026 2440
rect 11241 2431 11299 2437
rect 11241 2428 11253 2431
rect 11020 2400 11253 2428
rect 11020 2388 11026 2400
rect 11241 2397 11253 2400
rect 11287 2397 11299 2431
rect 11241 2391 11299 2397
rect 10318 2252 10324 2304
rect 10376 2292 10382 2304
rect 10505 2295 10563 2301
rect 10505 2292 10517 2295
rect 10376 2264 10517 2292
rect 10376 2252 10382 2264
rect 10505 2261 10517 2264
rect 10551 2261 10563 2295
rect 10505 2255 10563 2261
rect 1104 2202 18860 2224
rect 1104 2150 3610 2202
rect 3662 2150 3674 2202
rect 3726 2150 3738 2202
rect 3790 2150 3802 2202
rect 3854 2150 3866 2202
rect 3918 2150 13610 2202
rect 13662 2150 13674 2202
rect 13726 2150 13738 2202
rect 13790 2150 13802 2202
rect 13854 2150 13866 2202
rect 13918 2150 18860 2202
rect 1104 2128 18860 2150
<< via1 >>
rect 3610 17382 3662 17434
rect 3674 17382 3726 17434
rect 3738 17382 3790 17434
rect 3802 17382 3854 17434
rect 3866 17382 3918 17434
rect 13610 17382 13662 17434
rect 13674 17382 13726 17434
rect 13738 17382 13790 17434
rect 13802 17382 13854 17434
rect 13866 17382 13918 17434
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 3610 16294 3662 16346
rect 3674 16294 3726 16346
rect 3738 16294 3790 16346
rect 3802 16294 3854 16346
rect 3866 16294 3918 16346
rect 13610 16294 13662 16346
rect 13674 16294 13726 16346
rect 13738 16294 13790 16346
rect 13802 16294 13854 16346
rect 13866 16294 13918 16346
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 3610 15206 3662 15258
rect 3674 15206 3726 15258
rect 3738 15206 3790 15258
rect 3802 15206 3854 15258
rect 3866 15206 3918 15258
rect 13610 15206 13662 15258
rect 13674 15206 13726 15258
rect 13738 15206 13790 15258
rect 13802 15206 13854 15258
rect 13866 15206 13918 15258
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 3610 14118 3662 14170
rect 3674 14118 3726 14170
rect 3738 14118 3790 14170
rect 3802 14118 3854 14170
rect 3866 14118 3918 14170
rect 13610 14118 13662 14170
rect 13674 14118 13726 14170
rect 13738 14118 13790 14170
rect 13802 14118 13854 14170
rect 13866 14118 13918 14170
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 3610 13030 3662 13082
rect 3674 13030 3726 13082
rect 3738 13030 3790 13082
rect 3802 13030 3854 13082
rect 3866 13030 3918 13082
rect 13610 13030 13662 13082
rect 13674 13030 13726 13082
rect 13738 13030 13790 13082
rect 13802 13030 13854 13082
rect 13866 13030 13918 13082
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 3610 11942 3662 11994
rect 3674 11942 3726 11994
rect 3738 11942 3790 11994
rect 3802 11942 3854 11994
rect 3866 11942 3918 11994
rect 13610 11942 13662 11994
rect 13674 11942 13726 11994
rect 13738 11942 13790 11994
rect 13802 11942 13854 11994
rect 13866 11942 13918 11994
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 3610 10854 3662 10906
rect 3674 10854 3726 10906
rect 3738 10854 3790 10906
rect 3802 10854 3854 10906
rect 3866 10854 3918 10906
rect 13610 10854 13662 10906
rect 13674 10854 13726 10906
rect 13738 10854 13790 10906
rect 13802 10854 13854 10906
rect 13866 10854 13918 10906
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 10692 10004 10744 10056
rect 18420 9911 18472 9920
rect 18420 9877 18429 9911
rect 18429 9877 18463 9911
rect 18463 9877 18472 9911
rect 18420 9868 18472 9877
rect 3610 9766 3662 9818
rect 3674 9766 3726 9818
rect 3738 9766 3790 9818
rect 3802 9766 3854 9818
rect 3866 9766 3918 9818
rect 13610 9766 13662 9818
rect 13674 9766 13726 9818
rect 13738 9766 13790 9818
rect 13802 9766 13854 9818
rect 13866 9766 13918 9818
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 3610 8678 3662 8730
rect 3674 8678 3726 8730
rect 3738 8678 3790 8730
rect 3802 8678 3854 8730
rect 3866 8678 3918 8730
rect 13610 8678 13662 8730
rect 13674 8678 13726 8730
rect 13738 8678 13790 8730
rect 13802 8678 13854 8730
rect 13866 8678 13918 8730
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 3610 7590 3662 7642
rect 3674 7590 3726 7642
rect 3738 7590 3790 7642
rect 3802 7590 3854 7642
rect 3866 7590 3918 7642
rect 13610 7590 13662 7642
rect 13674 7590 13726 7642
rect 13738 7590 13790 7642
rect 13802 7590 13854 7642
rect 13866 7590 13918 7642
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 3610 6502 3662 6554
rect 3674 6502 3726 6554
rect 3738 6502 3790 6554
rect 3802 6502 3854 6554
rect 3866 6502 3918 6554
rect 13610 6502 13662 6554
rect 13674 6502 13726 6554
rect 13738 6502 13790 6554
rect 13802 6502 13854 6554
rect 13866 6502 13918 6554
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 3610 5414 3662 5466
rect 3674 5414 3726 5466
rect 3738 5414 3790 5466
rect 3802 5414 3854 5466
rect 3866 5414 3918 5466
rect 13610 5414 13662 5466
rect 13674 5414 13726 5466
rect 13738 5414 13790 5466
rect 13802 5414 13854 5466
rect 13866 5414 13918 5466
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 3610 4326 3662 4378
rect 3674 4326 3726 4378
rect 3738 4326 3790 4378
rect 3802 4326 3854 4378
rect 3866 4326 3918 4378
rect 13610 4326 13662 4378
rect 13674 4326 13726 4378
rect 13738 4326 13790 4378
rect 13802 4326 13854 4378
rect 13866 4326 13918 4378
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 10692 3655 10744 3664
rect 10692 3621 10701 3655
rect 10701 3621 10735 3655
rect 10735 3621 10744 3655
rect 10692 3612 10744 3621
rect 10232 3587 10284 3596
rect 10232 3553 10241 3587
rect 10241 3553 10275 3587
rect 10275 3553 10284 3587
rect 10232 3544 10284 3553
rect 10048 3476 10100 3528
rect 3610 3238 3662 3290
rect 3674 3238 3726 3290
rect 3738 3238 3790 3290
rect 3802 3238 3854 3290
rect 3866 3238 3918 3290
rect 13610 3238 13662 3290
rect 13674 3238 13726 3290
rect 13738 3238 13790 3290
rect 13802 3238 13854 3290
rect 13866 3238 13918 3290
rect 10232 3179 10284 3188
rect 10232 3145 10241 3179
rect 10241 3145 10275 3179
rect 10275 3145 10284 3179
rect 10232 3136 10284 3145
rect 10324 3043 10376 3052
rect 10324 3009 10333 3043
rect 10333 3009 10367 3043
rect 10367 3009 10376 3043
rect 10324 3000 10376 3009
rect 9956 2975 10008 2984
rect 9956 2941 9965 2975
rect 9965 2941 9999 2975
rect 9999 2941 10008 2975
rect 9956 2932 10008 2941
rect 11060 2864 11112 2916
rect 10692 2796 10744 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 10048 2592 10100 2644
rect 10324 2592 10376 2644
rect 11060 2635 11112 2644
rect 11060 2601 11069 2635
rect 11069 2601 11103 2635
rect 11103 2601 11112 2635
rect 11060 2592 11112 2601
rect 9956 2567 10008 2576
rect 9956 2533 9965 2567
rect 9965 2533 9999 2567
rect 9999 2533 10008 2567
rect 9956 2524 10008 2533
rect 9036 2388 9088 2440
rect 9680 2388 9732 2440
rect 10048 2431 10100 2440
rect 10048 2397 10057 2431
rect 10057 2397 10091 2431
rect 10091 2397 10100 2431
rect 10048 2388 10100 2397
rect 10692 2431 10744 2440
rect 10692 2397 10701 2431
rect 10701 2397 10735 2431
rect 10735 2397 10744 2431
rect 10692 2388 10744 2397
rect 10968 2388 11020 2440
rect 10324 2252 10376 2304
rect 3610 2150 3662 2202
rect 3674 2150 3726 2202
rect 3738 2150 3790 2202
rect 3802 2150 3854 2202
rect 3866 2150 3918 2202
rect 13610 2150 13662 2202
rect 13674 2150 13726 2202
rect 13738 2150 13790 2202
rect 13802 2150 13854 2202
rect 13866 2150 13918 2202
<< metal2 >>
rect 3610 17436 3918 17445
rect 3610 17434 3616 17436
rect 3672 17434 3696 17436
rect 3752 17434 3776 17436
rect 3832 17434 3856 17436
rect 3912 17434 3918 17436
rect 3672 17382 3674 17434
rect 3854 17382 3856 17434
rect 3610 17380 3616 17382
rect 3672 17380 3696 17382
rect 3752 17380 3776 17382
rect 3832 17380 3856 17382
rect 3912 17380 3918 17382
rect 3610 17371 3918 17380
rect 13610 17436 13918 17445
rect 13610 17434 13616 17436
rect 13672 17434 13696 17436
rect 13752 17434 13776 17436
rect 13832 17434 13856 17436
rect 13912 17434 13918 17436
rect 13672 17382 13674 17434
rect 13854 17382 13856 17434
rect 13610 17380 13616 17382
rect 13672 17380 13696 17382
rect 13752 17380 13776 17382
rect 13832 17380 13856 17382
rect 13912 17380 13918 17382
rect 13610 17371 13918 17380
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 3610 16348 3918 16357
rect 3610 16346 3616 16348
rect 3672 16346 3696 16348
rect 3752 16346 3776 16348
rect 3832 16346 3856 16348
rect 3912 16346 3918 16348
rect 3672 16294 3674 16346
rect 3854 16294 3856 16346
rect 3610 16292 3616 16294
rect 3672 16292 3696 16294
rect 3752 16292 3776 16294
rect 3832 16292 3856 16294
rect 3912 16292 3918 16294
rect 3610 16283 3918 16292
rect 13610 16348 13918 16357
rect 13610 16346 13616 16348
rect 13672 16346 13696 16348
rect 13752 16346 13776 16348
rect 13832 16346 13856 16348
rect 13912 16346 13918 16348
rect 13672 16294 13674 16346
rect 13854 16294 13856 16346
rect 13610 16292 13616 16294
rect 13672 16292 13696 16294
rect 13752 16292 13776 16294
rect 13832 16292 13856 16294
rect 13912 16292 13918 16294
rect 13610 16283 13918 16292
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 3610 15260 3918 15269
rect 3610 15258 3616 15260
rect 3672 15258 3696 15260
rect 3752 15258 3776 15260
rect 3832 15258 3856 15260
rect 3912 15258 3918 15260
rect 3672 15206 3674 15258
rect 3854 15206 3856 15258
rect 3610 15204 3616 15206
rect 3672 15204 3696 15206
rect 3752 15204 3776 15206
rect 3832 15204 3856 15206
rect 3912 15204 3918 15206
rect 3610 15195 3918 15204
rect 13610 15260 13918 15269
rect 13610 15258 13616 15260
rect 13672 15258 13696 15260
rect 13752 15258 13776 15260
rect 13832 15258 13856 15260
rect 13912 15258 13918 15260
rect 13672 15206 13674 15258
rect 13854 15206 13856 15258
rect 13610 15204 13616 15206
rect 13672 15204 13696 15206
rect 13752 15204 13776 15206
rect 13832 15204 13856 15206
rect 13912 15204 13918 15206
rect 13610 15195 13918 15204
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 3610 14172 3918 14181
rect 3610 14170 3616 14172
rect 3672 14170 3696 14172
rect 3752 14170 3776 14172
rect 3832 14170 3856 14172
rect 3912 14170 3918 14172
rect 3672 14118 3674 14170
rect 3854 14118 3856 14170
rect 3610 14116 3616 14118
rect 3672 14116 3696 14118
rect 3752 14116 3776 14118
rect 3832 14116 3856 14118
rect 3912 14116 3918 14118
rect 3610 14107 3918 14116
rect 13610 14172 13918 14181
rect 13610 14170 13616 14172
rect 13672 14170 13696 14172
rect 13752 14170 13776 14172
rect 13832 14170 13856 14172
rect 13912 14170 13918 14172
rect 13672 14118 13674 14170
rect 13854 14118 13856 14170
rect 13610 14116 13616 14118
rect 13672 14116 13696 14118
rect 13752 14116 13776 14118
rect 13832 14116 13856 14118
rect 13912 14116 13918 14118
rect 13610 14107 13918 14116
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 3610 13084 3918 13093
rect 3610 13082 3616 13084
rect 3672 13082 3696 13084
rect 3752 13082 3776 13084
rect 3832 13082 3856 13084
rect 3912 13082 3918 13084
rect 3672 13030 3674 13082
rect 3854 13030 3856 13082
rect 3610 13028 3616 13030
rect 3672 13028 3696 13030
rect 3752 13028 3776 13030
rect 3832 13028 3856 13030
rect 3912 13028 3918 13030
rect 3610 13019 3918 13028
rect 13610 13084 13918 13093
rect 13610 13082 13616 13084
rect 13672 13082 13696 13084
rect 13752 13082 13776 13084
rect 13832 13082 13856 13084
rect 13912 13082 13918 13084
rect 13672 13030 13674 13082
rect 13854 13030 13856 13082
rect 13610 13028 13616 13030
rect 13672 13028 13696 13030
rect 13752 13028 13776 13030
rect 13832 13028 13856 13030
rect 13912 13028 13918 13030
rect 13610 13019 13918 13028
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 3610 11996 3918 12005
rect 3610 11994 3616 11996
rect 3672 11994 3696 11996
rect 3752 11994 3776 11996
rect 3832 11994 3856 11996
rect 3912 11994 3918 11996
rect 3672 11942 3674 11994
rect 3854 11942 3856 11994
rect 3610 11940 3616 11942
rect 3672 11940 3696 11942
rect 3752 11940 3776 11942
rect 3832 11940 3856 11942
rect 3912 11940 3918 11942
rect 3610 11931 3918 11940
rect 13610 11996 13918 12005
rect 13610 11994 13616 11996
rect 13672 11994 13696 11996
rect 13752 11994 13776 11996
rect 13832 11994 13856 11996
rect 13912 11994 13918 11996
rect 13672 11942 13674 11994
rect 13854 11942 13856 11994
rect 13610 11940 13616 11942
rect 13672 11940 13696 11942
rect 13752 11940 13776 11942
rect 13832 11940 13856 11942
rect 13912 11940 13918 11942
rect 13610 11931 13918 11940
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 3610 10908 3918 10917
rect 3610 10906 3616 10908
rect 3672 10906 3696 10908
rect 3752 10906 3776 10908
rect 3832 10906 3856 10908
rect 3912 10906 3918 10908
rect 3672 10854 3674 10906
rect 3854 10854 3856 10906
rect 3610 10852 3616 10854
rect 3672 10852 3696 10854
rect 3752 10852 3776 10854
rect 3832 10852 3856 10854
rect 3912 10852 3918 10854
rect 3610 10843 3918 10852
rect 13610 10908 13918 10917
rect 13610 10906 13616 10908
rect 13672 10906 13696 10908
rect 13752 10906 13776 10908
rect 13832 10906 13856 10908
rect 13912 10906 13918 10908
rect 13672 10854 13674 10906
rect 13854 10854 13856 10906
rect 13610 10852 13616 10854
rect 13672 10852 13696 10854
rect 13752 10852 13776 10854
rect 13832 10852 13856 10854
rect 13912 10852 13918 10854
rect 13610 10843 13918 10852
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 3610 9820 3918 9829
rect 3610 9818 3616 9820
rect 3672 9818 3696 9820
rect 3752 9818 3776 9820
rect 3832 9818 3856 9820
rect 3912 9818 3918 9820
rect 3672 9766 3674 9818
rect 3854 9766 3856 9818
rect 3610 9764 3616 9766
rect 3672 9764 3696 9766
rect 3752 9764 3776 9766
rect 3832 9764 3856 9766
rect 3912 9764 3918 9766
rect 3610 9755 3918 9764
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 3610 8732 3918 8741
rect 3610 8730 3616 8732
rect 3672 8730 3696 8732
rect 3752 8730 3776 8732
rect 3832 8730 3856 8732
rect 3912 8730 3918 8732
rect 3672 8678 3674 8730
rect 3854 8678 3856 8730
rect 3610 8676 3616 8678
rect 3672 8676 3696 8678
rect 3752 8676 3776 8678
rect 3832 8676 3856 8678
rect 3912 8676 3918 8678
rect 3610 8667 3918 8676
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 3610 7644 3918 7653
rect 3610 7642 3616 7644
rect 3672 7642 3696 7644
rect 3752 7642 3776 7644
rect 3832 7642 3856 7644
rect 3912 7642 3918 7644
rect 3672 7590 3674 7642
rect 3854 7590 3856 7642
rect 3610 7588 3616 7590
rect 3672 7588 3696 7590
rect 3752 7588 3776 7590
rect 3832 7588 3856 7590
rect 3912 7588 3918 7590
rect 3610 7579 3918 7588
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 3610 6556 3918 6565
rect 3610 6554 3616 6556
rect 3672 6554 3696 6556
rect 3752 6554 3776 6556
rect 3832 6554 3856 6556
rect 3912 6554 3918 6556
rect 3672 6502 3674 6554
rect 3854 6502 3856 6554
rect 3610 6500 3616 6502
rect 3672 6500 3696 6502
rect 3752 6500 3776 6502
rect 3832 6500 3856 6502
rect 3912 6500 3918 6502
rect 3610 6491 3918 6500
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 3610 5468 3918 5477
rect 3610 5466 3616 5468
rect 3672 5466 3696 5468
rect 3752 5466 3776 5468
rect 3832 5466 3856 5468
rect 3912 5466 3918 5468
rect 3672 5414 3674 5466
rect 3854 5414 3856 5466
rect 3610 5412 3616 5414
rect 3672 5412 3696 5414
rect 3752 5412 3776 5414
rect 3832 5412 3856 5414
rect 3912 5412 3918 5414
rect 3610 5403 3918 5412
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 3610 4380 3918 4389
rect 3610 4378 3616 4380
rect 3672 4378 3696 4380
rect 3752 4378 3776 4380
rect 3832 4378 3856 4380
rect 3912 4378 3918 4380
rect 3672 4326 3674 4378
rect 3854 4326 3856 4378
rect 3610 4324 3616 4326
rect 3672 4324 3696 4326
rect 3752 4324 3776 4326
rect 3832 4324 3856 4326
rect 3912 4324 3918 4326
rect 3610 4315 3918 4324
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 10704 3670 10732 9998
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 13610 9820 13918 9829
rect 13610 9818 13616 9820
rect 13672 9818 13696 9820
rect 13752 9818 13776 9820
rect 13832 9818 13856 9820
rect 13912 9818 13918 9820
rect 13672 9766 13674 9818
rect 13854 9766 13856 9818
rect 13610 9764 13616 9766
rect 13672 9764 13696 9766
rect 13752 9764 13776 9766
rect 13832 9764 13856 9766
rect 13912 9764 13918 9766
rect 13610 9755 13918 9764
rect 18432 9625 18460 9862
rect 18418 9616 18474 9625
rect 18418 9551 18474 9560
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 13610 8732 13918 8741
rect 13610 8730 13616 8732
rect 13672 8730 13696 8732
rect 13752 8730 13776 8732
rect 13832 8730 13856 8732
rect 13912 8730 13918 8732
rect 13672 8678 13674 8730
rect 13854 8678 13856 8730
rect 13610 8676 13616 8678
rect 13672 8676 13696 8678
rect 13752 8676 13776 8678
rect 13832 8676 13856 8678
rect 13912 8676 13918 8678
rect 13610 8667 13918 8676
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 13610 7644 13918 7653
rect 13610 7642 13616 7644
rect 13672 7642 13696 7644
rect 13752 7642 13776 7644
rect 13832 7642 13856 7644
rect 13912 7642 13918 7644
rect 13672 7590 13674 7642
rect 13854 7590 13856 7642
rect 13610 7588 13616 7590
rect 13672 7588 13696 7590
rect 13752 7588 13776 7590
rect 13832 7588 13856 7590
rect 13912 7588 13918 7590
rect 13610 7579 13918 7588
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 13610 6556 13918 6565
rect 13610 6554 13616 6556
rect 13672 6554 13696 6556
rect 13752 6554 13776 6556
rect 13832 6554 13856 6556
rect 13912 6554 13918 6556
rect 13672 6502 13674 6554
rect 13854 6502 13856 6554
rect 13610 6500 13616 6502
rect 13672 6500 13696 6502
rect 13752 6500 13776 6502
rect 13832 6500 13856 6502
rect 13912 6500 13918 6502
rect 13610 6491 13918 6500
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 13610 5468 13918 5477
rect 13610 5466 13616 5468
rect 13672 5466 13696 5468
rect 13752 5466 13776 5468
rect 13832 5466 13856 5468
rect 13912 5466 13918 5468
rect 13672 5414 13674 5466
rect 13854 5414 13856 5466
rect 13610 5412 13616 5414
rect 13672 5412 13696 5414
rect 13752 5412 13776 5414
rect 13832 5412 13856 5414
rect 13912 5412 13918 5414
rect 13610 5403 13918 5412
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 13610 4380 13918 4389
rect 13610 4378 13616 4380
rect 13672 4378 13696 4380
rect 13752 4378 13776 4380
rect 13832 4378 13856 4380
rect 13912 4378 13918 4380
rect 13672 4326 13674 4378
rect 13854 4326 13856 4378
rect 13610 4324 13616 4326
rect 13672 4324 13696 4326
rect 13752 4324 13776 4326
rect 13832 4324 13856 4326
rect 13912 4324 13918 4326
rect 13610 4315 13918 4324
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 3610 3292 3918 3301
rect 3610 3290 3616 3292
rect 3672 3290 3696 3292
rect 3752 3290 3776 3292
rect 3832 3290 3856 3292
rect 3912 3290 3918 3292
rect 3672 3238 3674 3290
rect 3854 3238 3856 3290
rect 3610 3236 3616 3238
rect 3672 3236 3696 3238
rect 3752 3236 3776 3238
rect 3832 3236 3856 3238
rect 3912 3236 3918 3238
rect 3610 3227 3918 3236
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 9968 2582 9996 2926
rect 10060 2650 10088 3470
rect 10244 3194 10272 3538
rect 13610 3292 13918 3301
rect 13610 3290 13616 3292
rect 13672 3290 13696 3292
rect 13752 3290 13776 3292
rect 13832 3290 13856 3292
rect 13912 3290 13918 3292
rect 13672 3238 13674 3290
rect 13854 3238 13856 3290
rect 13610 3236 13616 3238
rect 13672 3236 13696 3238
rect 13752 3236 13776 3238
rect 13832 3236 13856 3238
rect 13912 3236 13918 3238
rect 13610 3227 13918 3236
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10336 2650 10364 2994
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 9956 2576 10008 2582
rect 9956 2518 10008 2524
rect 10060 2446 10088 2586
rect 10704 2446 10732 2790
rect 11072 2650 11100 2858
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 3610 2204 3918 2213
rect 3610 2202 3616 2204
rect 3672 2202 3696 2204
rect 3752 2202 3776 2204
rect 3832 2202 3856 2204
rect 3912 2202 3918 2204
rect 3672 2150 3674 2202
rect 3854 2150 3856 2202
rect 3610 2148 3616 2150
rect 3672 2148 3696 2150
rect 3752 2148 3776 2150
rect 3832 2148 3856 2150
rect 3912 2148 3918 2150
rect 3610 2139 3918 2148
rect 9048 800 9076 2382
rect 9692 800 9720 2382
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 10336 800 10364 2246
rect 10980 800 11008 2382
rect 13610 2204 13918 2213
rect 13610 2202 13616 2204
rect 13672 2202 13696 2204
rect 13752 2202 13776 2204
rect 13832 2202 13856 2204
rect 13912 2202 13918 2204
rect 13672 2150 13674 2202
rect 13854 2150 13856 2202
rect 13610 2148 13616 2150
rect 13672 2148 13696 2150
rect 13752 2148 13776 2150
rect 13832 2148 13856 2150
rect 13912 2148 13918 2150
rect 13610 2139 13918 2148
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
<< via2 >>
rect 3616 17434 3672 17436
rect 3696 17434 3752 17436
rect 3776 17434 3832 17436
rect 3856 17434 3912 17436
rect 3616 17382 3662 17434
rect 3662 17382 3672 17434
rect 3696 17382 3726 17434
rect 3726 17382 3738 17434
rect 3738 17382 3752 17434
rect 3776 17382 3790 17434
rect 3790 17382 3802 17434
rect 3802 17382 3832 17434
rect 3856 17382 3866 17434
rect 3866 17382 3912 17434
rect 3616 17380 3672 17382
rect 3696 17380 3752 17382
rect 3776 17380 3832 17382
rect 3856 17380 3912 17382
rect 13616 17434 13672 17436
rect 13696 17434 13752 17436
rect 13776 17434 13832 17436
rect 13856 17434 13912 17436
rect 13616 17382 13662 17434
rect 13662 17382 13672 17434
rect 13696 17382 13726 17434
rect 13726 17382 13738 17434
rect 13738 17382 13752 17434
rect 13776 17382 13790 17434
rect 13790 17382 13802 17434
rect 13802 17382 13832 17434
rect 13856 17382 13866 17434
rect 13866 17382 13912 17434
rect 13616 17380 13672 17382
rect 13696 17380 13752 17382
rect 13776 17380 13832 17382
rect 13856 17380 13912 17382
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 3616 16346 3672 16348
rect 3696 16346 3752 16348
rect 3776 16346 3832 16348
rect 3856 16346 3912 16348
rect 3616 16294 3662 16346
rect 3662 16294 3672 16346
rect 3696 16294 3726 16346
rect 3726 16294 3738 16346
rect 3738 16294 3752 16346
rect 3776 16294 3790 16346
rect 3790 16294 3802 16346
rect 3802 16294 3832 16346
rect 3856 16294 3866 16346
rect 3866 16294 3912 16346
rect 3616 16292 3672 16294
rect 3696 16292 3752 16294
rect 3776 16292 3832 16294
rect 3856 16292 3912 16294
rect 13616 16346 13672 16348
rect 13696 16346 13752 16348
rect 13776 16346 13832 16348
rect 13856 16346 13912 16348
rect 13616 16294 13662 16346
rect 13662 16294 13672 16346
rect 13696 16294 13726 16346
rect 13726 16294 13738 16346
rect 13738 16294 13752 16346
rect 13776 16294 13790 16346
rect 13790 16294 13802 16346
rect 13802 16294 13832 16346
rect 13856 16294 13866 16346
rect 13866 16294 13912 16346
rect 13616 16292 13672 16294
rect 13696 16292 13752 16294
rect 13776 16292 13832 16294
rect 13856 16292 13912 16294
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 3616 15258 3672 15260
rect 3696 15258 3752 15260
rect 3776 15258 3832 15260
rect 3856 15258 3912 15260
rect 3616 15206 3662 15258
rect 3662 15206 3672 15258
rect 3696 15206 3726 15258
rect 3726 15206 3738 15258
rect 3738 15206 3752 15258
rect 3776 15206 3790 15258
rect 3790 15206 3802 15258
rect 3802 15206 3832 15258
rect 3856 15206 3866 15258
rect 3866 15206 3912 15258
rect 3616 15204 3672 15206
rect 3696 15204 3752 15206
rect 3776 15204 3832 15206
rect 3856 15204 3912 15206
rect 13616 15258 13672 15260
rect 13696 15258 13752 15260
rect 13776 15258 13832 15260
rect 13856 15258 13912 15260
rect 13616 15206 13662 15258
rect 13662 15206 13672 15258
rect 13696 15206 13726 15258
rect 13726 15206 13738 15258
rect 13738 15206 13752 15258
rect 13776 15206 13790 15258
rect 13790 15206 13802 15258
rect 13802 15206 13832 15258
rect 13856 15206 13866 15258
rect 13866 15206 13912 15258
rect 13616 15204 13672 15206
rect 13696 15204 13752 15206
rect 13776 15204 13832 15206
rect 13856 15204 13912 15206
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 3616 14170 3672 14172
rect 3696 14170 3752 14172
rect 3776 14170 3832 14172
rect 3856 14170 3912 14172
rect 3616 14118 3662 14170
rect 3662 14118 3672 14170
rect 3696 14118 3726 14170
rect 3726 14118 3738 14170
rect 3738 14118 3752 14170
rect 3776 14118 3790 14170
rect 3790 14118 3802 14170
rect 3802 14118 3832 14170
rect 3856 14118 3866 14170
rect 3866 14118 3912 14170
rect 3616 14116 3672 14118
rect 3696 14116 3752 14118
rect 3776 14116 3832 14118
rect 3856 14116 3912 14118
rect 13616 14170 13672 14172
rect 13696 14170 13752 14172
rect 13776 14170 13832 14172
rect 13856 14170 13912 14172
rect 13616 14118 13662 14170
rect 13662 14118 13672 14170
rect 13696 14118 13726 14170
rect 13726 14118 13738 14170
rect 13738 14118 13752 14170
rect 13776 14118 13790 14170
rect 13790 14118 13802 14170
rect 13802 14118 13832 14170
rect 13856 14118 13866 14170
rect 13866 14118 13912 14170
rect 13616 14116 13672 14118
rect 13696 14116 13752 14118
rect 13776 14116 13832 14118
rect 13856 14116 13912 14118
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 3616 13082 3672 13084
rect 3696 13082 3752 13084
rect 3776 13082 3832 13084
rect 3856 13082 3912 13084
rect 3616 13030 3662 13082
rect 3662 13030 3672 13082
rect 3696 13030 3726 13082
rect 3726 13030 3738 13082
rect 3738 13030 3752 13082
rect 3776 13030 3790 13082
rect 3790 13030 3802 13082
rect 3802 13030 3832 13082
rect 3856 13030 3866 13082
rect 3866 13030 3912 13082
rect 3616 13028 3672 13030
rect 3696 13028 3752 13030
rect 3776 13028 3832 13030
rect 3856 13028 3912 13030
rect 13616 13082 13672 13084
rect 13696 13082 13752 13084
rect 13776 13082 13832 13084
rect 13856 13082 13912 13084
rect 13616 13030 13662 13082
rect 13662 13030 13672 13082
rect 13696 13030 13726 13082
rect 13726 13030 13738 13082
rect 13738 13030 13752 13082
rect 13776 13030 13790 13082
rect 13790 13030 13802 13082
rect 13802 13030 13832 13082
rect 13856 13030 13866 13082
rect 13866 13030 13912 13082
rect 13616 13028 13672 13030
rect 13696 13028 13752 13030
rect 13776 13028 13832 13030
rect 13856 13028 13912 13030
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 3616 11994 3672 11996
rect 3696 11994 3752 11996
rect 3776 11994 3832 11996
rect 3856 11994 3912 11996
rect 3616 11942 3662 11994
rect 3662 11942 3672 11994
rect 3696 11942 3726 11994
rect 3726 11942 3738 11994
rect 3738 11942 3752 11994
rect 3776 11942 3790 11994
rect 3790 11942 3802 11994
rect 3802 11942 3832 11994
rect 3856 11942 3866 11994
rect 3866 11942 3912 11994
rect 3616 11940 3672 11942
rect 3696 11940 3752 11942
rect 3776 11940 3832 11942
rect 3856 11940 3912 11942
rect 13616 11994 13672 11996
rect 13696 11994 13752 11996
rect 13776 11994 13832 11996
rect 13856 11994 13912 11996
rect 13616 11942 13662 11994
rect 13662 11942 13672 11994
rect 13696 11942 13726 11994
rect 13726 11942 13738 11994
rect 13738 11942 13752 11994
rect 13776 11942 13790 11994
rect 13790 11942 13802 11994
rect 13802 11942 13832 11994
rect 13856 11942 13866 11994
rect 13866 11942 13912 11994
rect 13616 11940 13672 11942
rect 13696 11940 13752 11942
rect 13776 11940 13832 11942
rect 13856 11940 13912 11942
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 3616 10906 3672 10908
rect 3696 10906 3752 10908
rect 3776 10906 3832 10908
rect 3856 10906 3912 10908
rect 3616 10854 3662 10906
rect 3662 10854 3672 10906
rect 3696 10854 3726 10906
rect 3726 10854 3738 10906
rect 3738 10854 3752 10906
rect 3776 10854 3790 10906
rect 3790 10854 3802 10906
rect 3802 10854 3832 10906
rect 3856 10854 3866 10906
rect 3866 10854 3912 10906
rect 3616 10852 3672 10854
rect 3696 10852 3752 10854
rect 3776 10852 3832 10854
rect 3856 10852 3912 10854
rect 13616 10906 13672 10908
rect 13696 10906 13752 10908
rect 13776 10906 13832 10908
rect 13856 10906 13912 10908
rect 13616 10854 13662 10906
rect 13662 10854 13672 10906
rect 13696 10854 13726 10906
rect 13726 10854 13738 10906
rect 13738 10854 13752 10906
rect 13776 10854 13790 10906
rect 13790 10854 13802 10906
rect 13802 10854 13832 10906
rect 13856 10854 13866 10906
rect 13866 10854 13912 10906
rect 13616 10852 13672 10854
rect 13696 10852 13752 10854
rect 13776 10852 13832 10854
rect 13856 10852 13912 10854
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 3616 9818 3672 9820
rect 3696 9818 3752 9820
rect 3776 9818 3832 9820
rect 3856 9818 3912 9820
rect 3616 9766 3662 9818
rect 3662 9766 3672 9818
rect 3696 9766 3726 9818
rect 3726 9766 3738 9818
rect 3738 9766 3752 9818
rect 3776 9766 3790 9818
rect 3790 9766 3802 9818
rect 3802 9766 3832 9818
rect 3856 9766 3866 9818
rect 3866 9766 3912 9818
rect 3616 9764 3672 9766
rect 3696 9764 3752 9766
rect 3776 9764 3832 9766
rect 3856 9764 3912 9766
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 3616 8730 3672 8732
rect 3696 8730 3752 8732
rect 3776 8730 3832 8732
rect 3856 8730 3912 8732
rect 3616 8678 3662 8730
rect 3662 8678 3672 8730
rect 3696 8678 3726 8730
rect 3726 8678 3738 8730
rect 3738 8678 3752 8730
rect 3776 8678 3790 8730
rect 3790 8678 3802 8730
rect 3802 8678 3832 8730
rect 3856 8678 3866 8730
rect 3866 8678 3912 8730
rect 3616 8676 3672 8678
rect 3696 8676 3752 8678
rect 3776 8676 3832 8678
rect 3856 8676 3912 8678
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 3616 7642 3672 7644
rect 3696 7642 3752 7644
rect 3776 7642 3832 7644
rect 3856 7642 3912 7644
rect 3616 7590 3662 7642
rect 3662 7590 3672 7642
rect 3696 7590 3726 7642
rect 3726 7590 3738 7642
rect 3738 7590 3752 7642
rect 3776 7590 3790 7642
rect 3790 7590 3802 7642
rect 3802 7590 3832 7642
rect 3856 7590 3866 7642
rect 3866 7590 3912 7642
rect 3616 7588 3672 7590
rect 3696 7588 3752 7590
rect 3776 7588 3832 7590
rect 3856 7588 3912 7590
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 3616 6554 3672 6556
rect 3696 6554 3752 6556
rect 3776 6554 3832 6556
rect 3856 6554 3912 6556
rect 3616 6502 3662 6554
rect 3662 6502 3672 6554
rect 3696 6502 3726 6554
rect 3726 6502 3738 6554
rect 3738 6502 3752 6554
rect 3776 6502 3790 6554
rect 3790 6502 3802 6554
rect 3802 6502 3832 6554
rect 3856 6502 3866 6554
rect 3866 6502 3912 6554
rect 3616 6500 3672 6502
rect 3696 6500 3752 6502
rect 3776 6500 3832 6502
rect 3856 6500 3912 6502
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 3616 5466 3672 5468
rect 3696 5466 3752 5468
rect 3776 5466 3832 5468
rect 3856 5466 3912 5468
rect 3616 5414 3662 5466
rect 3662 5414 3672 5466
rect 3696 5414 3726 5466
rect 3726 5414 3738 5466
rect 3738 5414 3752 5466
rect 3776 5414 3790 5466
rect 3790 5414 3802 5466
rect 3802 5414 3832 5466
rect 3856 5414 3866 5466
rect 3866 5414 3912 5466
rect 3616 5412 3672 5414
rect 3696 5412 3752 5414
rect 3776 5412 3832 5414
rect 3856 5412 3912 5414
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 3616 4378 3672 4380
rect 3696 4378 3752 4380
rect 3776 4378 3832 4380
rect 3856 4378 3912 4380
rect 3616 4326 3662 4378
rect 3662 4326 3672 4378
rect 3696 4326 3726 4378
rect 3726 4326 3738 4378
rect 3738 4326 3752 4378
rect 3776 4326 3790 4378
rect 3790 4326 3802 4378
rect 3802 4326 3832 4378
rect 3856 4326 3866 4378
rect 3866 4326 3912 4378
rect 3616 4324 3672 4326
rect 3696 4324 3752 4326
rect 3776 4324 3832 4326
rect 3856 4324 3912 4326
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 13616 9818 13672 9820
rect 13696 9818 13752 9820
rect 13776 9818 13832 9820
rect 13856 9818 13912 9820
rect 13616 9766 13662 9818
rect 13662 9766 13672 9818
rect 13696 9766 13726 9818
rect 13726 9766 13738 9818
rect 13738 9766 13752 9818
rect 13776 9766 13790 9818
rect 13790 9766 13802 9818
rect 13802 9766 13832 9818
rect 13856 9766 13866 9818
rect 13866 9766 13912 9818
rect 13616 9764 13672 9766
rect 13696 9764 13752 9766
rect 13776 9764 13832 9766
rect 13856 9764 13912 9766
rect 18418 9560 18474 9616
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 13616 8730 13672 8732
rect 13696 8730 13752 8732
rect 13776 8730 13832 8732
rect 13856 8730 13912 8732
rect 13616 8678 13662 8730
rect 13662 8678 13672 8730
rect 13696 8678 13726 8730
rect 13726 8678 13738 8730
rect 13738 8678 13752 8730
rect 13776 8678 13790 8730
rect 13790 8678 13802 8730
rect 13802 8678 13832 8730
rect 13856 8678 13866 8730
rect 13866 8678 13912 8730
rect 13616 8676 13672 8678
rect 13696 8676 13752 8678
rect 13776 8676 13832 8678
rect 13856 8676 13912 8678
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 13616 7642 13672 7644
rect 13696 7642 13752 7644
rect 13776 7642 13832 7644
rect 13856 7642 13912 7644
rect 13616 7590 13662 7642
rect 13662 7590 13672 7642
rect 13696 7590 13726 7642
rect 13726 7590 13738 7642
rect 13738 7590 13752 7642
rect 13776 7590 13790 7642
rect 13790 7590 13802 7642
rect 13802 7590 13832 7642
rect 13856 7590 13866 7642
rect 13866 7590 13912 7642
rect 13616 7588 13672 7590
rect 13696 7588 13752 7590
rect 13776 7588 13832 7590
rect 13856 7588 13912 7590
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 13616 6554 13672 6556
rect 13696 6554 13752 6556
rect 13776 6554 13832 6556
rect 13856 6554 13912 6556
rect 13616 6502 13662 6554
rect 13662 6502 13672 6554
rect 13696 6502 13726 6554
rect 13726 6502 13738 6554
rect 13738 6502 13752 6554
rect 13776 6502 13790 6554
rect 13790 6502 13802 6554
rect 13802 6502 13832 6554
rect 13856 6502 13866 6554
rect 13866 6502 13912 6554
rect 13616 6500 13672 6502
rect 13696 6500 13752 6502
rect 13776 6500 13832 6502
rect 13856 6500 13912 6502
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 13616 5466 13672 5468
rect 13696 5466 13752 5468
rect 13776 5466 13832 5468
rect 13856 5466 13912 5468
rect 13616 5414 13662 5466
rect 13662 5414 13672 5466
rect 13696 5414 13726 5466
rect 13726 5414 13738 5466
rect 13738 5414 13752 5466
rect 13776 5414 13790 5466
rect 13790 5414 13802 5466
rect 13802 5414 13832 5466
rect 13856 5414 13866 5466
rect 13866 5414 13912 5466
rect 13616 5412 13672 5414
rect 13696 5412 13752 5414
rect 13776 5412 13832 5414
rect 13856 5412 13912 5414
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 13616 4378 13672 4380
rect 13696 4378 13752 4380
rect 13776 4378 13832 4380
rect 13856 4378 13912 4380
rect 13616 4326 13662 4378
rect 13662 4326 13672 4378
rect 13696 4326 13726 4378
rect 13726 4326 13738 4378
rect 13738 4326 13752 4378
rect 13776 4326 13790 4378
rect 13790 4326 13802 4378
rect 13802 4326 13832 4378
rect 13856 4326 13866 4378
rect 13866 4326 13912 4378
rect 13616 4324 13672 4326
rect 13696 4324 13752 4326
rect 13776 4324 13832 4326
rect 13856 4324 13912 4326
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 3616 3290 3672 3292
rect 3696 3290 3752 3292
rect 3776 3290 3832 3292
rect 3856 3290 3912 3292
rect 3616 3238 3662 3290
rect 3662 3238 3672 3290
rect 3696 3238 3726 3290
rect 3726 3238 3738 3290
rect 3738 3238 3752 3290
rect 3776 3238 3790 3290
rect 3790 3238 3802 3290
rect 3802 3238 3832 3290
rect 3856 3238 3866 3290
rect 3866 3238 3912 3290
rect 3616 3236 3672 3238
rect 3696 3236 3752 3238
rect 3776 3236 3832 3238
rect 3856 3236 3912 3238
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 13616 3290 13672 3292
rect 13696 3290 13752 3292
rect 13776 3290 13832 3292
rect 13856 3290 13912 3292
rect 13616 3238 13662 3290
rect 13662 3238 13672 3290
rect 13696 3238 13726 3290
rect 13726 3238 13738 3290
rect 13738 3238 13752 3290
rect 13776 3238 13790 3290
rect 13790 3238 13802 3290
rect 13802 3238 13832 3290
rect 13856 3238 13866 3290
rect 13866 3238 13912 3290
rect 13616 3236 13672 3238
rect 13696 3236 13752 3238
rect 13776 3236 13832 3238
rect 13856 3236 13912 3238
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 3616 2202 3672 2204
rect 3696 2202 3752 2204
rect 3776 2202 3832 2204
rect 3856 2202 3912 2204
rect 3616 2150 3662 2202
rect 3662 2150 3672 2202
rect 3696 2150 3726 2202
rect 3726 2150 3738 2202
rect 3738 2150 3752 2202
rect 3776 2150 3790 2202
rect 3790 2150 3802 2202
rect 3802 2150 3832 2202
rect 3856 2150 3866 2202
rect 3866 2150 3912 2202
rect 3616 2148 3672 2150
rect 3696 2148 3752 2150
rect 3776 2148 3832 2150
rect 3856 2148 3912 2150
rect 13616 2202 13672 2204
rect 13696 2202 13752 2204
rect 13776 2202 13832 2204
rect 13856 2202 13912 2204
rect 13616 2150 13662 2202
rect 13662 2150 13672 2202
rect 13696 2150 13726 2202
rect 13726 2150 13738 2202
rect 13738 2150 13752 2202
rect 13776 2150 13790 2202
rect 13790 2150 13802 2202
rect 13802 2150 13832 2202
rect 13856 2150 13866 2202
rect 13866 2150 13912 2202
rect 13616 2148 13672 2150
rect 13696 2148 13752 2150
rect 13776 2148 13832 2150
rect 13856 2148 13912 2150
<< metal3 >>
rect 3606 17440 3922 17441
rect 3606 17376 3612 17440
rect 3676 17376 3692 17440
rect 3756 17376 3772 17440
rect 3836 17376 3852 17440
rect 3916 17376 3922 17440
rect 3606 17375 3922 17376
rect 13606 17440 13922 17441
rect 13606 17376 13612 17440
rect 13676 17376 13692 17440
rect 13756 17376 13772 17440
rect 13836 17376 13852 17440
rect 13916 17376 13922 17440
rect 13606 17375 13922 17376
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 3606 16352 3922 16353
rect 3606 16288 3612 16352
rect 3676 16288 3692 16352
rect 3756 16288 3772 16352
rect 3836 16288 3852 16352
rect 3916 16288 3922 16352
rect 3606 16287 3922 16288
rect 13606 16352 13922 16353
rect 13606 16288 13612 16352
rect 13676 16288 13692 16352
rect 13756 16288 13772 16352
rect 13836 16288 13852 16352
rect 13916 16288 13922 16352
rect 13606 16287 13922 16288
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 3606 15264 3922 15265
rect 3606 15200 3612 15264
rect 3676 15200 3692 15264
rect 3756 15200 3772 15264
rect 3836 15200 3852 15264
rect 3916 15200 3922 15264
rect 3606 15199 3922 15200
rect 13606 15264 13922 15265
rect 13606 15200 13612 15264
rect 13676 15200 13692 15264
rect 13756 15200 13772 15264
rect 13836 15200 13852 15264
rect 13916 15200 13922 15264
rect 13606 15199 13922 15200
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 3606 14176 3922 14177
rect 3606 14112 3612 14176
rect 3676 14112 3692 14176
rect 3756 14112 3772 14176
rect 3836 14112 3852 14176
rect 3916 14112 3922 14176
rect 3606 14111 3922 14112
rect 13606 14176 13922 14177
rect 13606 14112 13612 14176
rect 13676 14112 13692 14176
rect 13756 14112 13772 14176
rect 13836 14112 13852 14176
rect 13916 14112 13922 14176
rect 13606 14111 13922 14112
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 3606 13088 3922 13089
rect 3606 13024 3612 13088
rect 3676 13024 3692 13088
rect 3756 13024 3772 13088
rect 3836 13024 3852 13088
rect 3916 13024 3922 13088
rect 3606 13023 3922 13024
rect 13606 13088 13922 13089
rect 13606 13024 13612 13088
rect 13676 13024 13692 13088
rect 13756 13024 13772 13088
rect 13836 13024 13852 13088
rect 13916 13024 13922 13088
rect 13606 13023 13922 13024
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 3606 12000 3922 12001
rect 3606 11936 3612 12000
rect 3676 11936 3692 12000
rect 3756 11936 3772 12000
rect 3836 11936 3852 12000
rect 3916 11936 3922 12000
rect 3606 11935 3922 11936
rect 13606 12000 13922 12001
rect 13606 11936 13612 12000
rect 13676 11936 13692 12000
rect 13756 11936 13772 12000
rect 13836 11936 13852 12000
rect 13916 11936 13922 12000
rect 13606 11935 13922 11936
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 3606 10912 3922 10913
rect 3606 10848 3612 10912
rect 3676 10848 3692 10912
rect 3756 10848 3772 10912
rect 3836 10848 3852 10912
rect 3916 10848 3922 10912
rect 3606 10847 3922 10848
rect 13606 10912 13922 10913
rect 13606 10848 13612 10912
rect 13676 10848 13692 10912
rect 13756 10848 13772 10912
rect 13836 10848 13852 10912
rect 13916 10848 13922 10912
rect 13606 10847 13922 10848
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 3606 9824 3922 9825
rect 3606 9760 3612 9824
rect 3676 9760 3692 9824
rect 3756 9760 3772 9824
rect 3836 9760 3852 9824
rect 3916 9760 3922 9824
rect 3606 9759 3922 9760
rect 13606 9824 13922 9825
rect 13606 9760 13612 9824
rect 13676 9760 13692 9824
rect 13756 9760 13772 9824
rect 13836 9760 13852 9824
rect 13916 9760 13922 9824
rect 13606 9759 13922 9760
rect 18413 9618 18479 9621
rect 19200 9618 20000 9648
rect 18413 9616 20000 9618
rect 18413 9560 18418 9616
rect 18474 9560 20000 9616
rect 18413 9558 20000 9560
rect 18413 9555 18479 9558
rect 19200 9528 20000 9558
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 3606 8736 3922 8737
rect 3606 8672 3612 8736
rect 3676 8672 3692 8736
rect 3756 8672 3772 8736
rect 3836 8672 3852 8736
rect 3916 8672 3922 8736
rect 3606 8671 3922 8672
rect 13606 8736 13922 8737
rect 13606 8672 13612 8736
rect 13676 8672 13692 8736
rect 13756 8672 13772 8736
rect 13836 8672 13852 8736
rect 13916 8672 13922 8736
rect 13606 8671 13922 8672
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 3606 7648 3922 7649
rect 3606 7584 3612 7648
rect 3676 7584 3692 7648
rect 3756 7584 3772 7648
rect 3836 7584 3852 7648
rect 3916 7584 3922 7648
rect 3606 7583 3922 7584
rect 13606 7648 13922 7649
rect 13606 7584 13612 7648
rect 13676 7584 13692 7648
rect 13756 7584 13772 7648
rect 13836 7584 13852 7648
rect 13916 7584 13922 7648
rect 13606 7583 13922 7584
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 3606 6560 3922 6561
rect 3606 6496 3612 6560
rect 3676 6496 3692 6560
rect 3756 6496 3772 6560
rect 3836 6496 3852 6560
rect 3916 6496 3922 6560
rect 3606 6495 3922 6496
rect 13606 6560 13922 6561
rect 13606 6496 13612 6560
rect 13676 6496 13692 6560
rect 13756 6496 13772 6560
rect 13836 6496 13852 6560
rect 13916 6496 13922 6560
rect 13606 6495 13922 6496
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 3606 5472 3922 5473
rect 3606 5408 3612 5472
rect 3676 5408 3692 5472
rect 3756 5408 3772 5472
rect 3836 5408 3852 5472
rect 3916 5408 3922 5472
rect 3606 5407 3922 5408
rect 13606 5472 13922 5473
rect 13606 5408 13612 5472
rect 13676 5408 13692 5472
rect 13756 5408 13772 5472
rect 13836 5408 13852 5472
rect 13916 5408 13922 5472
rect 13606 5407 13922 5408
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 3606 4384 3922 4385
rect 3606 4320 3612 4384
rect 3676 4320 3692 4384
rect 3756 4320 3772 4384
rect 3836 4320 3852 4384
rect 3916 4320 3922 4384
rect 3606 4319 3922 4320
rect 13606 4384 13922 4385
rect 13606 4320 13612 4384
rect 13676 4320 13692 4384
rect 13756 4320 13772 4384
rect 13836 4320 13852 4384
rect 13916 4320 13922 4384
rect 13606 4319 13922 4320
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 3606 3296 3922 3297
rect 3606 3232 3612 3296
rect 3676 3232 3692 3296
rect 3756 3232 3772 3296
rect 3836 3232 3852 3296
rect 3916 3232 3922 3296
rect 3606 3231 3922 3232
rect 13606 3296 13922 3297
rect 13606 3232 13612 3296
rect 13676 3232 13692 3296
rect 13756 3232 13772 3296
rect 13836 3232 13852 3296
rect 13916 3232 13922 3296
rect 13606 3231 13922 3232
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 3606 2208 3922 2209
rect 3606 2144 3612 2208
rect 3676 2144 3692 2208
rect 3756 2144 3772 2208
rect 3836 2144 3852 2208
rect 3916 2144 3922 2208
rect 3606 2143 3922 2144
rect 13606 2208 13922 2209
rect 13606 2144 13612 2208
rect 13676 2144 13692 2208
rect 13756 2144 13772 2208
rect 13836 2144 13852 2208
rect 13916 2144 13922 2208
rect 13606 2143 13922 2144
<< via3 >>
rect 3612 17436 3676 17440
rect 3612 17380 3616 17436
rect 3616 17380 3672 17436
rect 3672 17380 3676 17436
rect 3612 17376 3676 17380
rect 3692 17436 3756 17440
rect 3692 17380 3696 17436
rect 3696 17380 3752 17436
rect 3752 17380 3756 17436
rect 3692 17376 3756 17380
rect 3772 17436 3836 17440
rect 3772 17380 3776 17436
rect 3776 17380 3832 17436
rect 3832 17380 3836 17436
rect 3772 17376 3836 17380
rect 3852 17436 3916 17440
rect 3852 17380 3856 17436
rect 3856 17380 3912 17436
rect 3912 17380 3916 17436
rect 3852 17376 3916 17380
rect 13612 17436 13676 17440
rect 13612 17380 13616 17436
rect 13616 17380 13672 17436
rect 13672 17380 13676 17436
rect 13612 17376 13676 17380
rect 13692 17436 13756 17440
rect 13692 17380 13696 17436
rect 13696 17380 13752 17436
rect 13752 17380 13756 17436
rect 13692 17376 13756 17380
rect 13772 17436 13836 17440
rect 13772 17380 13776 17436
rect 13776 17380 13832 17436
rect 13832 17380 13836 17436
rect 13772 17376 13836 17380
rect 13852 17436 13916 17440
rect 13852 17380 13856 17436
rect 13856 17380 13912 17436
rect 13912 17380 13916 17436
rect 13852 17376 13916 17380
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 3612 16348 3676 16352
rect 3612 16292 3616 16348
rect 3616 16292 3672 16348
rect 3672 16292 3676 16348
rect 3612 16288 3676 16292
rect 3692 16348 3756 16352
rect 3692 16292 3696 16348
rect 3696 16292 3752 16348
rect 3752 16292 3756 16348
rect 3692 16288 3756 16292
rect 3772 16348 3836 16352
rect 3772 16292 3776 16348
rect 3776 16292 3832 16348
rect 3832 16292 3836 16348
rect 3772 16288 3836 16292
rect 3852 16348 3916 16352
rect 3852 16292 3856 16348
rect 3856 16292 3912 16348
rect 3912 16292 3916 16348
rect 3852 16288 3916 16292
rect 13612 16348 13676 16352
rect 13612 16292 13616 16348
rect 13616 16292 13672 16348
rect 13672 16292 13676 16348
rect 13612 16288 13676 16292
rect 13692 16348 13756 16352
rect 13692 16292 13696 16348
rect 13696 16292 13752 16348
rect 13752 16292 13756 16348
rect 13692 16288 13756 16292
rect 13772 16348 13836 16352
rect 13772 16292 13776 16348
rect 13776 16292 13832 16348
rect 13832 16292 13836 16348
rect 13772 16288 13836 16292
rect 13852 16348 13916 16352
rect 13852 16292 13856 16348
rect 13856 16292 13912 16348
rect 13912 16292 13916 16348
rect 13852 16288 13916 16292
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 3612 15260 3676 15264
rect 3612 15204 3616 15260
rect 3616 15204 3672 15260
rect 3672 15204 3676 15260
rect 3612 15200 3676 15204
rect 3692 15260 3756 15264
rect 3692 15204 3696 15260
rect 3696 15204 3752 15260
rect 3752 15204 3756 15260
rect 3692 15200 3756 15204
rect 3772 15260 3836 15264
rect 3772 15204 3776 15260
rect 3776 15204 3832 15260
rect 3832 15204 3836 15260
rect 3772 15200 3836 15204
rect 3852 15260 3916 15264
rect 3852 15204 3856 15260
rect 3856 15204 3912 15260
rect 3912 15204 3916 15260
rect 3852 15200 3916 15204
rect 13612 15260 13676 15264
rect 13612 15204 13616 15260
rect 13616 15204 13672 15260
rect 13672 15204 13676 15260
rect 13612 15200 13676 15204
rect 13692 15260 13756 15264
rect 13692 15204 13696 15260
rect 13696 15204 13752 15260
rect 13752 15204 13756 15260
rect 13692 15200 13756 15204
rect 13772 15260 13836 15264
rect 13772 15204 13776 15260
rect 13776 15204 13832 15260
rect 13832 15204 13836 15260
rect 13772 15200 13836 15204
rect 13852 15260 13916 15264
rect 13852 15204 13856 15260
rect 13856 15204 13912 15260
rect 13912 15204 13916 15260
rect 13852 15200 13916 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 3612 14172 3676 14176
rect 3612 14116 3616 14172
rect 3616 14116 3672 14172
rect 3672 14116 3676 14172
rect 3612 14112 3676 14116
rect 3692 14172 3756 14176
rect 3692 14116 3696 14172
rect 3696 14116 3752 14172
rect 3752 14116 3756 14172
rect 3692 14112 3756 14116
rect 3772 14172 3836 14176
rect 3772 14116 3776 14172
rect 3776 14116 3832 14172
rect 3832 14116 3836 14172
rect 3772 14112 3836 14116
rect 3852 14172 3916 14176
rect 3852 14116 3856 14172
rect 3856 14116 3912 14172
rect 3912 14116 3916 14172
rect 3852 14112 3916 14116
rect 13612 14172 13676 14176
rect 13612 14116 13616 14172
rect 13616 14116 13672 14172
rect 13672 14116 13676 14172
rect 13612 14112 13676 14116
rect 13692 14172 13756 14176
rect 13692 14116 13696 14172
rect 13696 14116 13752 14172
rect 13752 14116 13756 14172
rect 13692 14112 13756 14116
rect 13772 14172 13836 14176
rect 13772 14116 13776 14172
rect 13776 14116 13832 14172
rect 13832 14116 13836 14172
rect 13772 14112 13836 14116
rect 13852 14172 13916 14176
rect 13852 14116 13856 14172
rect 13856 14116 13912 14172
rect 13912 14116 13916 14172
rect 13852 14112 13916 14116
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 3612 13084 3676 13088
rect 3612 13028 3616 13084
rect 3616 13028 3672 13084
rect 3672 13028 3676 13084
rect 3612 13024 3676 13028
rect 3692 13084 3756 13088
rect 3692 13028 3696 13084
rect 3696 13028 3752 13084
rect 3752 13028 3756 13084
rect 3692 13024 3756 13028
rect 3772 13084 3836 13088
rect 3772 13028 3776 13084
rect 3776 13028 3832 13084
rect 3832 13028 3836 13084
rect 3772 13024 3836 13028
rect 3852 13084 3916 13088
rect 3852 13028 3856 13084
rect 3856 13028 3912 13084
rect 3912 13028 3916 13084
rect 3852 13024 3916 13028
rect 13612 13084 13676 13088
rect 13612 13028 13616 13084
rect 13616 13028 13672 13084
rect 13672 13028 13676 13084
rect 13612 13024 13676 13028
rect 13692 13084 13756 13088
rect 13692 13028 13696 13084
rect 13696 13028 13752 13084
rect 13752 13028 13756 13084
rect 13692 13024 13756 13028
rect 13772 13084 13836 13088
rect 13772 13028 13776 13084
rect 13776 13028 13832 13084
rect 13832 13028 13836 13084
rect 13772 13024 13836 13028
rect 13852 13084 13916 13088
rect 13852 13028 13856 13084
rect 13856 13028 13912 13084
rect 13912 13028 13916 13084
rect 13852 13024 13916 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 3612 11996 3676 12000
rect 3612 11940 3616 11996
rect 3616 11940 3672 11996
rect 3672 11940 3676 11996
rect 3612 11936 3676 11940
rect 3692 11996 3756 12000
rect 3692 11940 3696 11996
rect 3696 11940 3752 11996
rect 3752 11940 3756 11996
rect 3692 11936 3756 11940
rect 3772 11996 3836 12000
rect 3772 11940 3776 11996
rect 3776 11940 3832 11996
rect 3832 11940 3836 11996
rect 3772 11936 3836 11940
rect 3852 11996 3916 12000
rect 3852 11940 3856 11996
rect 3856 11940 3912 11996
rect 3912 11940 3916 11996
rect 3852 11936 3916 11940
rect 13612 11996 13676 12000
rect 13612 11940 13616 11996
rect 13616 11940 13672 11996
rect 13672 11940 13676 11996
rect 13612 11936 13676 11940
rect 13692 11996 13756 12000
rect 13692 11940 13696 11996
rect 13696 11940 13752 11996
rect 13752 11940 13756 11996
rect 13692 11936 13756 11940
rect 13772 11996 13836 12000
rect 13772 11940 13776 11996
rect 13776 11940 13832 11996
rect 13832 11940 13836 11996
rect 13772 11936 13836 11940
rect 13852 11996 13916 12000
rect 13852 11940 13856 11996
rect 13856 11940 13912 11996
rect 13912 11940 13916 11996
rect 13852 11936 13916 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 3612 10908 3676 10912
rect 3612 10852 3616 10908
rect 3616 10852 3672 10908
rect 3672 10852 3676 10908
rect 3612 10848 3676 10852
rect 3692 10908 3756 10912
rect 3692 10852 3696 10908
rect 3696 10852 3752 10908
rect 3752 10852 3756 10908
rect 3692 10848 3756 10852
rect 3772 10908 3836 10912
rect 3772 10852 3776 10908
rect 3776 10852 3832 10908
rect 3832 10852 3836 10908
rect 3772 10848 3836 10852
rect 3852 10908 3916 10912
rect 3852 10852 3856 10908
rect 3856 10852 3912 10908
rect 3912 10852 3916 10908
rect 3852 10848 3916 10852
rect 13612 10908 13676 10912
rect 13612 10852 13616 10908
rect 13616 10852 13672 10908
rect 13672 10852 13676 10908
rect 13612 10848 13676 10852
rect 13692 10908 13756 10912
rect 13692 10852 13696 10908
rect 13696 10852 13752 10908
rect 13752 10852 13756 10908
rect 13692 10848 13756 10852
rect 13772 10908 13836 10912
rect 13772 10852 13776 10908
rect 13776 10852 13832 10908
rect 13832 10852 13836 10908
rect 13772 10848 13836 10852
rect 13852 10908 13916 10912
rect 13852 10852 13856 10908
rect 13856 10852 13912 10908
rect 13912 10852 13916 10908
rect 13852 10848 13916 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 3612 9820 3676 9824
rect 3612 9764 3616 9820
rect 3616 9764 3672 9820
rect 3672 9764 3676 9820
rect 3612 9760 3676 9764
rect 3692 9820 3756 9824
rect 3692 9764 3696 9820
rect 3696 9764 3752 9820
rect 3752 9764 3756 9820
rect 3692 9760 3756 9764
rect 3772 9820 3836 9824
rect 3772 9764 3776 9820
rect 3776 9764 3832 9820
rect 3832 9764 3836 9820
rect 3772 9760 3836 9764
rect 3852 9820 3916 9824
rect 3852 9764 3856 9820
rect 3856 9764 3912 9820
rect 3912 9764 3916 9820
rect 3852 9760 3916 9764
rect 13612 9820 13676 9824
rect 13612 9764 13616 9820
rect 13616 9764 13672 9820
rect 13672 9764 13676 9820
rect 13612 9760 13676 9764
rect 13692 9820 13756 9824
rect 13692 9764 13696 9820
rect 13696 9764 13752 9820
rect 13752 9764 13756 9820
rect 13692 9760 13756 9764
rect 13772 9820 13836 9824
rect 13772 9764 13776 9820
rect 13776 9764 13832 9820
rect 13832 9764 13836 9820
rect 13772 9760 13836 9764
rect 13852 9820 13916 9824
rect 13852 9764 13856 9820
rect 13856 9764 13912 9820
rect 13912 9764 13916 9820
rect 13852 9760 13916 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 3612 8732 3676 8736
rect 3612 8676 3616 8732
rect 3616 8676 3672 8732
rect 3672 8676 3676 8732
rect 3612 8672 3676 8676
rect 3692 8732 3756 8736
rect 3692 8676 3696 8732
rect 3696 8676 3752 8732
rect 3752 8676 3756 8732
rect 3692 8672 3756 8676
rect 3772 8732 3836 8736
rect 3772 8676 3776 8732
rect 3776 8676 3832 8732
rect 3832 8676 3836 8732
rect 3772 8672 3836 8676
rect 3852 8732 3916 8736
rect 3852 8676 3856 8732
rect 3856 8676 3912 8732
rect 3912 8676 3916 8732
rect 3852 8672 3916 8676
rect 13612 8732 13676 8736
rect 13612 8676 13616 8732
rect 13616 8676 13672 8732
rect 13672 8676 13676 8732
rect 13612 8672 13676 8676
rect 13692 8732 13756 8736
rect 13692 8676 13696 8732
rect 13696 8676 13752 8732
rect 13752 8676 13756 8732
rect 13692 8672 13756 8676
rect 13772 8732 13836 8736
rect 13772 8676 13776 8732
rect 13776 8676 13832 8732
rect 13832 8676 13836 8732
rect 13772 8672 13836 8676
rect 13852 8732 13916 8736
rect 13852 8676 13856 8732
rect 13856 8676 13912 8732
rect 13912 8676 13916 8732
rect 13852 8672 13916 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 3612 7644 3676 7648
rect 3612 7588 3616 7644
rect 3616 7588 3672 7644
rect 3672 7588 3676 7644
rect 3612 7584 3676 7588
rect 3692 7644 3756 7648
rect 3692 7588 3696 7644
rect 3696 7588 3752 7644
rect 3752 7588 3756 7644
rect 3692 7584 3756 7588
rect 3772 7644 3836 7648
rect 3772 7588 3776 7644
rect 3776 7588 3832 7644
rect 3832 7588 3836 7644
rect 3772 7584 3836 7588
rect 3852 7644 3916 7648
rect 3852 7588 3856 7644
rect 3856 7588 3912 7644
rect 3912 7588 3916 7644
rect 3852 7584 3916 7588
rect 13612 7644 13676 7648
rect 13612 7588 13616 7644
rect 13616 7588 13672 7644
rect 13672 7588 13676 7644
rect 13612 7584 13676 7588
rect 13692 7644 13756 7648
rect 13692 7588 13696 7644
rect 13696 7588 13752 7644
rect 13752 7588 13756 7644
rect 13692 7584 13756 7588
rect 13772 7644 13836 7648
rect 13772 7588 13776 7644
rect 13776 7588 13832 7644
rect 13832 7588 13836 7644
rect 13772 7584 13836 7588
rect 13852 7644 13916 7648
rect 13852 7588 13856 7644
rect 13856 7588 13912 7644
rect 13912 7588 13916 7644
rect 13852 7584 13916 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 3612 6556 3676 6560
rect 3612 6500 3616 6556
rect 3616 6500 3672 6556
rect 3672 6500 3676 6556
rect 3612 6496 3676 6500
rect 3692 6556 3756 6560
rect 3692 6500 3696 6556
rect 3696 6500 3752 6556
rect 3752 6500 3756 6556
rect 3692 6496 3756 6500
rect 3772 6556 3836 6560
rect 3772 6500 3776 6556
rect 3776 6500 3832 6556
rect 3832 6500 3836 6556
rect 3772 6496 3836 6500
rect 3852 6556 3916 6560
rect 3852 6500 3856 6556
rect 3856 6500 3912 6556
rect 3912 6500 3916 6556
rect 3852 6496 3916 6500
rect 13612 6556 13676 6560
rect 13612 6500 13616 6556
rect 13616 6500 13672 6556
rect 13672 6500 13676 6556
rect 13612 6496 13676 6500
rect 13692 6556 13756 6560
rect 13692 6500 13696 6556
rect 13696 6500 13752 6556
rect 13752 6500 13756 6556
rect 13692 6496 13756 6500
rect 13772 6556 13836 6560
rect 13772 6500 13776 6556
rect 13776 6500 13832 6556
rect 13832 6500 13836 6556
rect 13772 6496 13836 6500
rect 13852 6556 13916 6560
rect 13852 6500 13856 6556
rect 13856 6500 13912 6556
rect 13912 6500 13916 6556
rect 13852 6496 13916 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 3612 5468 3676 5472
rect 3612 5412 3616 5468
rect 3616 5412 3672 5468
rect 3672 5412 3676 5468
rect 3612 5408 3676 5412
rect 3692 5468 3756 5472
rect 3692 5412 3696 5468
rect 3696 5412 3752 5468
rect 3752 5412 3756 5468
rect 3692 5408 3756 5412
rect 3772 5468 3836 5472
rect 3772 5412 3776 5468
rect 3776 5412 3832 5468
rect 3832 5412 3836 5468
rect 3772 5408 3836 5412
rect 3852 5468 3916 5472
rect 3852 5412 3856 5468
rect 3856 5412 3912 5468
rect 3912 5412 3916 5468
rect 3852 5408 3916 5412
rect 13612 5468 13676 5472
rect 13612 5412 13616 5468
rect 13616 5412 13672 5468
rect 13672 5412 13676 5468
rect 13612 5408 13676 5412
rect 13692 5468 13756 5472
rect 13692 5412 13696 5468
rect 13696 5412 13752 5468
rect 13752 5412 13756 5468
rect 13692 5408 13756 5412
rect 13772 5468 13836 5472
rect 13772 5412 13776 5468
rect 13776 5412 13832 5468
rect 13832 5412 13836 5468
rect 13772 5408 13836 5412
rect 13852 5468 13916 5472
rect 13852 5412 13856 5468
rect 13856 5412 13912 5468
rect 13912 5412 13916 5468
rect 13852 5408 13916 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 3612 4380 3676 4384
rect 3612 4324 3616 4380
rect 3616 4324 3672 4380
rect 3672 4324 3676 4380
rect 3612 4320 3676 4324
rect 3692 4380 3756 4384
rect 3692 4324 3696 4380
rect 3696 4324 3752 4380
rect 3752 4324 3756 4380
rect 3692 4320 3756 4324
rect 3772 4380 3836 4384
rect 3772 4324 3776 4380
rect 3776 4324 3832 4380
rect 3832 4324 3836 4380
rect 3772 4320 3836 4324
rect 3852 4380 3916 4384
rect 3852 4324 3856 4380
rect 3856 4324 3912 4380
rect 3912 4324 3916 4380
rect 3852 4320 3916 4324
rect 13612 4380 13676 4384
rect 13612 4324 13616 4380
rect 13616 4324 13672 4380
rect 13672 4324 13676 4380
rect 13612 4320 13676 4324
rect 13692 4380 13756 4384
rect 13692 4324 13696 4380
rect 13696 4324 13752 4380
rect 13752 4324 13756 4380
rect 13692 4320 13756 4324
rect 13772 4380 13836 4384
rect 13772 4324 13776 4380
rect 13776 4324 13832 4380
rect 13832 4324 13836 4380
rect 13772 4320 13836 4324
rect 13852 4380 13916 4384
rect 13852 4324 13856 4380
rect 13856 4324 13912 4380
rect 13912 4324 13916 4380
rect 13852 4320 13916 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 3612 3292 3676 3296
rect 3612 3236 3616 3292
rect 3616 3236 3672 3292
rect 3672 3236 3676 3292
rect 3612 3232 3676 3236
rect 3692 3292 3756 3296
rect 3692 3236 3696 3292
rect 3696 3236 3752 3292
rect 3752 3236 3756 3292
rect 3692 3232 3756 3236
rect 3772 3292 3836 3296
rect 3772 3236 3776 3292
rect 3776 3236 3832 3292
rect 3832 3236 3836 3292
rect 3772 3232 3836 3236
rect 3852 3292 3916 3296
rect 3852 3236 3856 3292
rect 3856 3236 3912 3292
rect 3912 3236 3916 3292
rect 3852 3232 3916 3236
rect 13612 3292 13676 3296
rect 13612 3236 13616 3292
rect 13616 3236 13672 3292
rect 13672 3236 13676 3292
rect 13612 3232 13676 3236
rect 13692 3292 13756 3296
rect 13692 3236 13696 3292
rect 13696 3236 13752 3292
rect 13752 3236 13756 3292
rect 13692 3232 13756 3236
rect 13772 3292 13836 3296
rect 13772 3236 13776 3292
rect 13776 3236 13832 3292
rect 13832 3236 13836 3292
rect 13772 3232 13836 3236
rect 13852 3292 13916 3296
rect 13852 3236 13856 3292
rect 13856 3236 13912 3292
rect 13912 3236 13916 3292
rect 13852 3232 13916 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 3612 2204 3676 2208
rect 3612 2148 3616 2204
rect 3616 2148 3672 2204
rect 3672 2148 3676 2204
rect 3612 2144 3676 2148
rect 3692 2204 3756 2208
rect 3692 2148 3696 2204
rect 3696 2148 3752 2204
rect 3752 2148 3756 2204
rect 3692 2144 3756 2148
rect 3772 2204 3836 2208
rect 3772 2148 3776 2204
rect 3776 2148 3832 2204
rect 3832 2148 3836 2204
rect 3772 2144 3836 2148
rect 3852 2204 3916 2208
rect 3852 2148 3856 2204
rect 3856 2148 3912 2204
rect 3912 2148 3916 2204
rect 3852 2144 3916 2148
rect 13612 2204 13676 2208
rect 13612 2148 13616 2204
rect 13616 2148 13672 2204
rect 13672 2148 13676 2204
rect 13612 2144 13676 2148
rect 13692 2204 13756 2208
rect 13692 2148 13696 2204
rect 13696 2148 13752 2204
rect 13752 2148 13756 2204
rect 13692 2144 13756 2148
rect 13772 2204 13836 2208
rect 13772 2148 13776 2204
rect 13776 2148 13832 2204
rect 13832 2148 13836 2204
rect 13772 2144 13836 2148
rect 13852 2204 13916 2208
rect 13852 2148 13856 2204
rect 13856 2148 13912 2204
rect 13912 2148 13916 2204
rect 13852 2144 13916 2148
<< metal4 >>
rect 2944 16896 3264 17456
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 14294 3264 14656
rect 2944 14058 2986 14294
rect 3222 14058 3264 14294
rect 2944 13632 3264 14058
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 4294 3264 4864
rect 2944 4058 2986 4294
rect 3222 4058 3264 4294
rect 2944 3840 3264 4058
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 3604 17440 3924 17456
rect 3604 17376 3612 17440
rect 3676 17376 3692 17440
rect 3756 17376 3772 17440
rect 3836 17376 3852 17440
rect 3916 17376 3924 17440
rect 3604 16352 3924 17376
rect 3604 16288 3612 16352
rect 3676 16288 3692 16352
rect 3756 16288 3772 16352
rect 3836 16288 3852 16352
rect 3916 16288 3924 16352
rect 3604 15264 3924 16288
rect 3604 15200 3612 15264
rect 3676 15200 3692 15264
rect 3756 15200 3772 15264
rect 3836 15200 3852 15264
rect 3916 15200 3924 15264
rect 3604 14954 3924 15200
rect 3604 14718 3646 14954
rect 3882 14718 3924 14954
rect 3604 14176 3924 14718
rect 3604 14112 3612 14176
rect 3676 14112 3692 14176
rect 3756 14112 3772 14176
rect 3836 14112 3852 14176
rect 3916 14112 3924 14176
rect 3604 13088 3924 14112
rect 3604 13024 3612 13088
rect 3676 13024 3692 13088
rect 3756 13024 3772 13088
rect 3836 13024 3852 13088
rect 3916 13024 3924 13088
rect 3604 12000 3924 13024
rect 3604 11936 3612 12000
rect 3676 11936 3692 12000
rect 3756 11936 3772 12000
rect 3836 11936 3852 12000
rect 3916 11936 3924 12000
rect 3604 10912 3924 11936
rect 3604 10848 3612 10912
rect 3676 10848 3692 10912
rect 3756 10848 3772 10912
rect 3836 10848 3852 10912
rect 3916 10848 3924 10912
rect 3604 9824 3924 10848
rect 3604 9760 3612 9824
rect 3676 9760 3692 9824
rect 3756 9760 3772 9824
rect 3836 9760 3852 9824
rect 3916 9760 3924 9824
rect 3604 8736 3924 9760
rect 3604 8672 3612 8736
rect 3676 8672 3692 8736
rect 3756 8672 3772 8736
rect 3836 8672 3852 8736
rect 3916 8672 3924 8736
rect 3604 7648 3924 8672
rect 3604 7584 3612 7648
rect 3676 7584 3692 7648
rect 3756 7584 3772 7648
rect 3836 7584 3852 7648
rect 3916 7584 3924 7648
rect 3604 6560 3924 7584
rect 3604 6496 3612 6560
rect 3676 6496 3692 6560
rect 3756 6496 3772 6560
rect 3836 6496 3852 6560
rect 3916 6496 3924 6560
rect 3604 5472 3924 6496
rect 3604 5408 3612 5472
rect 3676 5408 3692 5472
rect 3756 5408 3772 5472
rect 3836 5408 3852 5472
rect 3916 5408 3924 5472
rect 3604 4954 3924 5408
rect 3604 4718 3646 4954
rect 3882 4718 3924 4954
rect 3604 4384 3924 4718
rect 3604 4320 3612 4384
rect 3676 4320 3692 4384
rect 3756 4320 3772 4384
rect 3836 4320 3852 4384
rect 3916 4320 3924 4384
rect 3604 3296 3924 4320
rect 3604 3232 3612 3296
rect 3676 3232 3692 3296
rect 3756 3232 3772 3296
rect 3836 3232 3852 3296
rect 3916 3232 3924 3296
rect 3604 2208 3924 3232
rect 3604 2144 3612 2208
rect 3676 2144 3692 2208
rect 3756 2144 3772 2208
rect 3836 2144 3852 2208
rect 3916 2144 3924 2208
rect 3604 2128 3924 2144
rect 12944 16896 13264 17456
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 14294 13264 14656
rect 12944 14058 12986 14294
rect 13222 14058 13264 14294
rect 12944 13632 13264 14058
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 4294 13264 4864
rect 12944 4058 12986 4294
rect 13222 4058 13264 4294
rect 12944 3840 13264 4058
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 13604 17440 13924 17456
rect 13604 17376 13612 17440
rect 13676 17376 13692 17440
rect 13756 17376 13772 17440
rect 13836 17376 13852 17440
rect 13916 17376 13924 17440
rect 13604 16352 13924 17376
rect 13604 16288 13612 16352
rect 13676 16288 13692 16352
rect 13756 16288 13772 16352
rect 13836 16288 13852 16352
rect 13916 16288 13924 16352
rect 13604 15264 13924 16288
rect 13604 15200 13612 15264
rect 13676 15200 13692 15264
rect 13756 15200 13772 15264
rect 13836 15200 13852 15264
rect 13916 15200 13924 15264
rect 13604 14954 13924 15200
rect 13604 14718 13646 14954
rect 13882 14718 13924 14954
rect 13604 14176 13924 14718
rect 13604 14112 13612 14176
rect 13676 14112 13692 14176
rect 13756 14112 13772 14176
rect 13836 14112 13852 14176
rect 13916 14112 13924 14176
rect 13604 13088 13924 14112
rect 13604 13024 13612 13088
rect 13676 13024 13692 13088
rect 13756 13024 13772 13088
rect 13836 13024 13852 13088
rect 13916 13024 13924 13088
rect 13604 12000 13924 13024
rect 13604 11936 13612 12000
rect 13676 11936 13692 12000
rect 13756 11936 13772 12000
rect 13836 11936 13852 12000
rect 13916 11936 13924 12000
rect 13604 10912 13924 11936
rect 13604 10848 13612 10912
rect 13676 10848 13692 10912
rect 13756 10848 13772 10912
rect 13836 10848 13852 10912
rect 13916 10848 13924 10912
rect 13604 9824 13924 10848
rect 13604 9760 13612 9824
rect 13676 9760 13692 9824
rect 13756 9760 13772 9824
rect 13836 9760 13852 9824
rect 13916 9760 13924 9824
rect 13604 8736 13924 9760
rect 13604 8672 13612 8736
rect 13676 8672 13692 8736
rect 13756 8672 13772 8736
rect 13836 8672 13852 8736
rect 13916 8672 13924 8736
rect 13604 7648 13924 8672
rect 13604 7584 13612 7648
rect 13676 7584 13692 7648
rect 13756 7584 13772 7648
rect 13836 7584 13852 7648
rect 13916 7584 13924 7648
rect 13604 6560 13924 7584
rect 13604 6496 13612 6560
rect 13676 6496 13692 6560
rect 13756 6496 13772 6560
rect 13836 6496 13852 6560
rect 13916 6496 13924 6560
rect 13604 5472 13924 6496
rect 13604 5408 13612 5472
rect 13676 5408 13692 5472
rect 13756 5408 13772 5472
rect 13836 5408 13852 5472
rect 13916 5408 13924 5472
rect 13604 4954 13924 5408
rect 13604 4718 13646 4954
rect 13882 4718 13924 4954
rect 13604 4384 13924 4718
rect 13604 4320 13612 4384
rect 13676 4320 13692 4384
rect 13756 4320 13772 4384
rect 13836 4320 13852 4384
rect 13916 4320 13924 4384
rect 13604 3296 13924 4320
rect 13604 3232 13612 3296
rect 13676 3232 13692 3296
rect 13756 3232 13772 3296
rect 13836 3232 13852 3296
rect 13916 3232 13924 3296
rect 13604 2208 13924 3232
rect 13604 2144 13612 2208
rect 13676 2144 13692 2208
rect 13756 2144 13772 2208
rect 13836 2144 13852 2208
rect 13916 2144 13924 2208
rect 13604 2128 13924 2144
<< via4 >>
rect 2986 14058 3222 14294
rect 2986 4058 3222 4294
rect 3646 14718 3882 14954
rect 3646 4718 3882 4954
rect 12986 14058 13222 14294
rect 12986 4058 13222 4294
rect 13646 14718 13882 14954
rect 13646 4718 13882 4954
<< metal5 >>
rect 1056 14954 18908 14996
rect 1056 14718 3646 14954
rect 3882 14718 13646 14954
rect 13882 14718 18908 14954
rect 1056 14676 18908 14718
rect 1056 14294 18908 14336
rect 1056 14058 2986 14294
rect 3222 14058 12986 14294
rect 13222 14058 18908 14294
rect 1056 14016 18908 14058
rect 1056 4954 18908 4996
rect 1056 4718 3646 4954
rect 3882 4718 13646 4954
rect 13882 4718 18908 4954
rect 1056 4676 18908 4718
rect 1056 4294 18908 4336
rect 1056 4058 2986 4294
rect 3222 4058 12986 4294
rect 13222 4058 18908 4294
rect 1056 4016 18908 4058
use sky130_fd_sc_hd__o21ai_1  _3_
timestamp 1
transform 1 0 10304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _4_
timestamp 1
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _5_
timestamp 1
transform 1 0 10672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _6_
timestamp 1
transform 1 0 9660 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _7_
timestamp 1
transform 1 0 10120 0 1 3264
box -38 -48 682 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100
timestamp 1
transform 1 0 10304 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_105
timestamp 1
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636968456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636968456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636968456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636968456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_181
timestamp 1
transform 1 0 17756 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_189
timestamp 1
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636968456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636968456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636968456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636968456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636968456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636968456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636968456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636968456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_181
timestamp 1
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_189
timestamp 1
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636968456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636968456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636968456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636968456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_97
timestamp 1
transform 1 0 10028 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_105
timestamp 1636968456
transform 1 0 10764 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_117
timestamp 1636968456
transform 1 0 11868 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_129
timestamp 1
transform 1 0 12972 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636968456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636968456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636968456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636968456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_189
timestamp 1
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636968456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636968456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636968456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636968456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636968456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636968456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636968456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636968456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636968456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636968456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636968456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_181
timestamp 1
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636968456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636968456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636968456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636968456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636968456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636968456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636968456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636968456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636968456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636968456
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636968456
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636968456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_189
timestamp 1
transform 1 0 18492 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636968456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636968456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636968456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636968456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636968456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636968456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636968456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636968456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636968456
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636968456
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636968456
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636968456
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636968456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_181
timestamp 1
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_189
timestamp 1
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636968456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636968456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636968456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636968456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636968456
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636968456
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636968456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636968456
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636968456
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1636968456
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636968456
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636968456
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636968456
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636968456
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_189
timestamp 1
transform 1 0 18492 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636968456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636968456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636968456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636968456
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636968456
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636968456
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636968456
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1636968456
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636968456
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636968456
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1636968456
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1636968456
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636968456
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_181
timestamp 1
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_189
timestamp 1
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636968456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636968456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636968456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636968456
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636968456
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636968456
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636968456
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1636968456
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1636968456
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1636968456
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636968456
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636968456
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636968456
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1636968456
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_189
timestamp 1
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636968456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636968456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636968456
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1636968456
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636968456
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636968456
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1636968456
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1636968456
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636968456
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1636968456
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1636968456
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1636968456
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636968456
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_181
timestamp 1
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_189
timestamp 1
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636968456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636968456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636968456
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636968456
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1636968456
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1636968456
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636968456
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1636968456
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1636968456
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1636968456
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1636968456
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1636968456
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1636968456
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1636968456
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636968456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636968456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1636968456
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1636968456
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636968456
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1636968456
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1636968456
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1636968456
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1636968456
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1636968456
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1636968456
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1636968456
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1636968456
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_181
timestamp 1
transform 1 0 17756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_189
timestamp 1
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636968456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636968456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636968456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636968456
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1636968456
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1636968456
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1636968456
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1636968456
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1636968456
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1636968456
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1636968456
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1636968456
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1636968456
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1636968456
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636968456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636968456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636968456
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1636968456
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1636968456
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1636968456
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1636968456
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1636968456
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1636968456
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1636968456
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1636968456
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1636968456
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1636968456
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_181
timestamp 1
transform 1 0 17756 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_189
timestamp 1
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636968456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636968456
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636968456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1636968456
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1636968456
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1636968456
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1636968456
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1636968456
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1636968456
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1636968456
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1636968456
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1636968456
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1636968456
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_177
timestamp 1
transform 1 0 17388 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_185
timestamp 1
transform 1 0 18124 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636968456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636968456
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636968456
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1636968456
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1636968456
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1636968456
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1636968456
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1636968456
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1636968456
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1636968456
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1636968456
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1636968456
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1636968456
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_181
timestamp 1
transform 1 0 17756 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_189
timestamp 1
transform 1 0 18492 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636968456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636968456
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636968456
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1636968456
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1636968456
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1636968456
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1636968456
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1636968456
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1636968456
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1636968456
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1636968456
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1636968456
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1636968456
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1636968456
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636968456
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1636968456
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1636968456
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1636968456
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636968456
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1636968456
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1636968456
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1636968456
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1636968456
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1636968456
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1636968456
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1636968456
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1636968456
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_181
timestamp 1
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp 1
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636968456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636968456
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636968456
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1636968456
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1636968456
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1636968456
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1636968456
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1636968456
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1636968456
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1636968456
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1636968456
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1636968456
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1636968456
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1636968456
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_189
timestamp 1
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636968456
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636968456
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1636968456
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1636968456
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636968456
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1636968456
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1636968456
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1636968456
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1636968456
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1636968456
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1636968456
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1636968456
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1636968456
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_181
timestamp 1
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 1
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636968456
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1636968456
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636968456
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1636968456
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1636968456
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1636968456
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1636968456
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1636968456
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1636968456
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1636968456
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1636968456
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1636968456
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1636968456
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1636968456
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_189
timestamp 1
transform 1 0 18492 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636968456
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636968456
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1636968456
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1636968456
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1636968456
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1636968456
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1636968456
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1636968456
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1636968456
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1636968456
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1636968456
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1636968456
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1636968456
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_181
timestamp 1
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp 1
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636968456
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636968456
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636968456
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1636968456
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1636968456
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1636968456
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1636968456
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1636968456
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1636968456
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1636968456
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1636968456
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1636968456
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1636968456
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1636968456
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_189
timestamp 1
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636968456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1636968456
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1636968456
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1636968456
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1636968456
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1636968456
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1636968456
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1636968456
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1636968456
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1636968456
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1636968456
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1636968456
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1636968456
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_181
timestamp 1
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_189
timestamp 1
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636968456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636968456
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636968456
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1636968456
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1636968456
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1636968456
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1636968456
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1636968456
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1636968456
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1636968456
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1636968456
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1636968456
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1636968456
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1636968456
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_189
timestamp 1
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1636968456
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1636968456
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1636968456
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1636968456
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1636968456
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1636968456
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1636968456
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1636968456
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1636968456
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1636968456
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1636968456
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1636968456
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1636968456
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_181
timestamp 1
transform 1 0 17756 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_189
timestamp 1
transform 1 0 18492 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636968456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636968456
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636968456
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1636968456
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1636968456
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1636968456
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1636968456
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1636968456
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1636968456
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1636968456
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1636968456
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1636968456
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1636968456
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1636968456
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_189
timestamp 1
transform 1 0 18492 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1636968456
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1636968456
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_29
timestamp 1636968456
transform 1 0 3772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_41
timestamp 1636968456
transform 1 0 4876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1636968456
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1636968456
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_81
timestamp 1
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_85
timestamp 1636968456
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_97
timestamp 1636968456
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1636968456
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1636968456
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_137
timestamp 1
transform 1 0 13708 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_141
timestamp 1636968456
transform 1 0 14076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_153
timestamp 1636968456
transform 1 0 15180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1636968456
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_181
timestamp 1
transform 1 0 17756 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_189
timestamp 1
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1
transform -1 0 11316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1
transform -1 0 10764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1
transform 1 0 18216 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_28
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_29
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_30
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_31
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_32
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_33
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_34
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_35
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_36
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_37
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_38
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_39
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_40
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_41
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_42
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_43
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_44
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_45
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_46
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_47
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_48
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_49
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_50
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_51
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_52
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_53
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_54
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_55
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_56
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_57
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_59
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_61
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_62
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_63
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_64
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_65
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_66
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_67
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_68
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_69
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_70
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_71
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_72
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_73
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_74
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_75
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_76
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_83
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_84
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_85
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_86
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_87
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_88
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_89
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_90
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_91
timestamp 1
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_92
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_93
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_94
timestamp 1
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_95
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_96
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_97
timestamp 1
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_98
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_99
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_100
timestamp 1
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_101
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_102
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_103
timestamp 1
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_104
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_105
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_106
timestamp 1
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_107
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_108
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_109
timestamp 1
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_110
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_111
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_112
timestamp 1
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_113
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_114
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_115
timestamp 1
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_116
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_117
timestamp 1
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_118
timestamp 1
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_119
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_120
timestamp 1
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_121
timestamp 1
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_122
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_123
timestamp 1
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_124
timestamp 1
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_125
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_126
timestamp 1
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_127
timestamp 1
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_128
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_129
timestamp 1
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_130
timestamp 1
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_131
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_132
timestamp 1
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_133
timestamp 1
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_134
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_135
timestamp 1
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_136
timestamp 1
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_137
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_138
timestamp 1
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_139
timestamp 1
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_140
timestamp 1
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_141
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_142
timestamp 1
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_143
timestamp 1
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_144
timestamp 1
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_145
timestamp 1
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
<< labels >>
flabel metal4 s 3604 2128 3924 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 13604 2128 13924 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 4676 18908 4996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 14676 18908 14996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 4016 18908 4336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 14016 18908 14336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 a_i
port 2 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 b_i
port 3 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 cin_i
port 4 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 cout_o
port 5 nsew signal output
flabel metal3 s 19200 9528 20000 9648 0 FreeSans 480 0 0 0 sum_o
port 6 nsew signal output
rlabel metal1 9982 17408 9982 17408 0 VGND
rlabel metal1 9982 16864 9982 16864 0 VPWR
rlabel metal1 10258 2618 10258 2618 0 _0_
rlabel metal1 10718 2958 10718 2958 0 _1_
rlabel metal2 10258 3366 10258 3366 0 _2_
rlabel metal2 9706 1588 9706 1588 0 a_i
rlabel metal2 10994 1588 10994 1588 0 b_i
rlabel metal2 9062 1588 9062 1588 0 cin_i
rlabel metal2 10350 1520 10350 1520 0 cout_o
rlabel metal1 10258 2958 10258 2958 0 net1
rlabel metal1 10902 2958 10902 2958 0 net2
rlabel metal2 10074 2958 10074 2958 0 net3
rlabel metal2 10718 2618 10718 2618 0 net4
rlabel metal2 10718 6834 10718 6834 0 net5
rlabel metal2 18446 9741 18446 9741 0 sum_o
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
